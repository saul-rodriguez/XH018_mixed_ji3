************************************************************************
* auCdl Netlist:
* 
* Library Name:  INV_HV
* Top Cell Name: inv_hv
* View Name:     schematic
* Netlisted on:  Feb  5 07:19:00 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE METER
.PARAM



************************************************************************
* Library Name: INV_HV
* Cell Name:    inv_hv
* View Name:    schematic
************************************************************************

.SUBCKT inv_hv GNDHV IN OUT VDDHV VSUB
*.PININFO GNDHV:B IN:B OUT:B VDDHV:B VSUB:B
MM0 OUT IN GNDHV VSUB NEDIA W=40u L=1.25u M=1.0 $LDD[NEDIA]
RR0 VDDHV OUT 9999.84 $SUB=VSUB $[RPP1K1_3] $W=10u $L=103.425u M=1
.ENDS

