* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : inv                                          *
* Netlisted  : Sun Feb  4 10:15:44 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3) nem ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pe3) pem pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ne3_CDNS_707059739800                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ne3_CDNS_707059739800 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 ne3 L=3.5e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=0
.ends ne3_CDNS_707059739800

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pe3_CDNS_707059739801                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pe3_CDNS_707059739801 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 2 3 1 1 pe3 L=3e-07 W=2e-06 AD=9.6e-13 AS=9.6e-13 PD=4.96e-06 PS=4.96e-06 $X=0 $Y=0 $dt=1
.ends pe3_CDNS_707059739801

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv IN OUT VD VS
** N=4 EP=4 FDC=3
X0 VS OUT IN ne3_CDNS_707059739800 $T=2000 2040 0 0 $X=1200 $Y=1640
X1 VD OUT IN pe3_CDNS_707059739801 $T=2025 5870 0 0 $X=515 $Y=4840
D0 VS VD p_dnw3 AREA=8.321e-12 PJ=1.209e-05 perimeter=1.209e-05 $X=1115 $Y=5440 $dt=2
.ends inv
