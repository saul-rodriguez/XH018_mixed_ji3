* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : counter_lvs                                  *
* Netlisted  : Sat Feb  3 17:36:07 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3i) nemi ndiff(D) p1trm(G) ndiff(S) pwitrm(B)
*.DEVTMPLT 1 MP(pe3i) pemi pdiff(D) p1trm(G) pdiff(S) dnwtrm(B)
*.DEVTMPLT 2 D(p_ddnwmv) p_ddnwmv bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 3 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX2 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=6
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=6e-07 AD=2.96727e-13 AS=2.88e-13 PD=1.69091e-06 PS=2.16e-06 $X=620 $Y=950 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=2.016e-13 AS=3.56073e-13 PD=1.512e-06 PS=2.02909e-06 $X=1590 $Y=830 $dt=0
M2 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=4.648e-13 AS=1.344e-13 PD=3.52e-06 PS=1.008e-06 $X=2480 $Y=1070 $dt=0
M3 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=5.39943e-13 AS=5.28e-13 PD=2.20442e-06 PS=3.16e-06 $X=620 $Y=2410 $dt=1
M4 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=7.16507e-13 PD=1.87971e-06 PS=2.92528e-06 $X=1640 $Y=2410 $dt=1
M5 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=8.6265e-13 AS=2.751e-13 PD=4.56971e-06 PS=1.87971e-06 $X=2480 $Y=2410 $dt=1
.ends BUJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX0                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX0 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=4
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.923e-13 AS=2.016e-13 PD=2.005e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.923e-13 PD=1.8e-06 PS=2.005e-06 $X=1735 $Y=1130 $dt=0
M2 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=9e-07 AD=5.7805e-13 AS=4.32e-13 PD=2.33911e-06 PS=2.76e-06 $X=620 $Y=2410 $dt=1
M3 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.12e-06 AD=5.376e-13 AS=7.1935e-13 PD=3.2e-06 PS=2.91089e-06 $X=1785 $Y=2410 $dt=1
.ends BUJI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX16                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX16 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=39
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=2400 $Y=660 $dt=0
M3 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=3290 $Y=660 $dt=0
M4 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=4180 $Y=660 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.4475e-13 AS=2.403e-13 PD=1.44e-06 PS=1.43e-06 $X=5070 $Y=660 $dt=0
M6 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.63267e-13 AS=2.4475e-13 PD=1.95905e-06 PS=1.44e-06 $X=5970 $Y=660 $dt=0
M7 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.26533e-13 PD=1.34e-06 PS=1.76095e-06 $X=6940 $Y=750 $dt=0
M8 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=7830 $Y=750 $dt=0
M9 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=8800 $Y=750 $dt=0
M10 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=9690 $Y=750 $dt=0
M11 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=10660 $Y=750 $dt=0
M12 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=11550 $Y=750 $dt=0
M13 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=12520 $Y=750 $dt=0
M14 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=13410 $Y=750 $dt=0
M15 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=14380 $Y=750 $dt=0
M16 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=2.16e-13 PD=2.56e-06 PS=1.34e-06 $X=15270 $Y=750 $dt=0
M17 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M18 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M19 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M20 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M21 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M22 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
M23 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4645 $Y=2410 $dt=1
M24 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=5485 $Y=2410 $dt=1
M25 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6035 $Y=2410 $dt=1
M26 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6875 $Y=2410 $dt=1
M27 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=7425 $Y=2410 $dt=1
M28 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8265 $Y=2410 $dt=1
M29 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8815 $Y=2410 $dt=1
M30 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=9655 $Y=2410 $dt=1
M31 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=10205 $Y=2410 $dt=1
M32 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=11045 $Y=2410 $dt=1
M33 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=11595 $Y=2410 $dt=1
M34 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=12435 $Y=2410 $dt=1
M35 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=12985 $Y=2410 $dt=1
M36 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=13825 $Y=2410 $dt=1
M37 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=14375 $Y=2410 $dt=1
M38 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=1.15229e-12 AS=2.54913e-13 PD=4.89506e-06 PS=1.86506e-06 $X=15215 $Y=2410 $dt=1
.ends BUJI3VX16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY1JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY1JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=8 EP=4 FDC=8
M0 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.591e-13 AS=2.016e-13 PD=2.13e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 6 8 gnd3i! gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.415e-13 AS=3.591e-13 PD=1.99e-06 PS=2.13e-06 $X=1590 $Y=1400 $dt=0
M2 gnd3i! 6 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=2.6662e-13 AS=2.016e-13 PD=1.28565e-06 PS=1.8e-06 $X=2860 $Y=660 $dt=0
M3 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.3165e-13 AS=5.6498e-13 PD=2.75e-06 PS=2.72435e-06 $X=4625 $Y=660 $dt=0
M4 vdd3i! A 8 vdd3i! pe3i L=3e-07 W=6.7e-07 AD=4.61962e-13 AS=3.3835e-13 PD=2.62468e-06 PS=2.35e-06 $X=645 $Y=2680 $dt=1
M5 6 8 vdd3i! vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.00088e-13 AS=2.89588e-13 PD=1.76778e-06 PS=1.64532e-06 $X=1590 $Y=2680 $dt=1
M6 vdd3i! 6 7 vdd3i! pe3i L=7.5e-07 W=4.2e-07 AD=2.78313e-13 AS=2.00088e-13 PD=1.17049e-06 PS=1.76778e-06 $X=3110 $Y=3400 $dt=1
M7 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.191e-13 AS=9.34337e-13 PD=3.84e-06 PS=3.92951e-06 $X=4650 $Y=2410 $dt=1
.ends DLY1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY2JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY2JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=12 EP=4 FDC=12
M0 gnd3i! A 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.577e-13 AS=2.016e-13 PD=1.79e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 8 10 gnd3i! gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.548e-13 AS=3.577e-13 PD=1.7e-06 PS=1.79e-06 $X=1990 $Y=660 $dt=0
M2 8 10 9 gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.548e-13 AS=2.016e-13 PD=1.7e-06 PS=1.8e-06 $X=1990 $Y=1360 $dt=0
M3 gnd3i! 9 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=3.42444e-13 AS=2.1e-13 PD=1.66718e-06 PS=1.62e-06 $X=3950 $Y=660 $dt=0
M4 6 9 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=2.10588e-13 AS=2.1e-13 PD=1.81778e-06 PS=1.62e-06 $X=3950 $Y=1360 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=7.25656e-13 PD=2.74e-06 PS=3.53282e-06 $X=6310 $Y=660 $dt=0
M6 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.42937e-13 AS=3.535e-13 PD=2.69375e-06 PS=2.41e-06 $X=645 $Y=3120 $dt=1
M7 12 10 9 vdd3i! pe3i L=7.4e-07 W=4.2e-07 AD=2.8095e-13 AS=2.0035e-13 PD=1.785e-06 PS=1.77071e-06 $X=2050 $Y=2640 $dt=1
M8 12 10 vdd3i! vdd3i! pe3i L=7.4e-07 W=4.2e-07 AD=2.8095e-13 AS=3.25762e-13 PD=1.785e-06 PS=1.61625e-06 $X=2050 $Y=3400 $dt=1
M9 6 9 11 vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.856e-13 AS=2.479e-13 PD=2.2e-06 PS=1.715e-06 $X=4030 $Y=2660 $dt=1
M10 vdd3i! 9 11 vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.62018e-13 AS=2.479e-13 PD=1.40689e-06 PS=1.715e-06 $X=4030 $Y=3400 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=8.79632e-13 PD=3.83e-06 PS=4.72311e-06 $X=6335 $Y=2410 $dt=1
.ends DLY2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=4
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.44533e-13 AS=2.016e-13 PD=1.44667e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=2.88e-13 AS=3.84267e-13 PD=2.28e-06 PS=2.27333e-06 $X=1590 $Y=890 $dt=0
M2 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=9e-07 AD=4.7931e-13 AS=4.32e-13 PD=1.95649e-06 PS=2.76e-06 $X=620 $Y=2410 $dt=1
M3 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=5.712e-13 AS=7.7739e-13 PD=3.70971e-06 PS=3.17322e-06 $X=1640 $Y=2410 $dt=1
.ends BUJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRQJI3VX2                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRQJI3VX2 vdd3i! gnd3i! D C Q
*.DEVICECLIMB
** N=20 EP=5 FDC=28
M0 gnd3i! 8 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=2.016e-13 PD=9.6e-07 PS=1.8e-06 $X=620 $Y=1000 $dt=0
M1 15 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=6.09e-14 AS=1.134e-13 PD=7.1e-07 PS=9.6e-07 $X=1510 $Y=1000 $dt=0
M2 8 12 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.30725e-13 AS=6.09e-14 PD=9.3e-07 PS=7.1e-07 $X=2150 $Y=1000 $dt=0
M3 14 13 8 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=2.17875e-13 PD=9.5e-07 PS=1.55e-06 $X=3040 $Y=960 $dt=0
M4 gnd3i! D 14 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=6.04277e-13 AS=8.75e-14 PD=3.74159e-06 PS=9.5e-07 $X=3640 $Y=960 $dt=0
M5 gnd3i! C 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.62566e-13 AS=2.016e-13 PD=2.24496e-06 PS=1.8e-06 $X=5070 $Y=1295 $dt=0
M6 12 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.62566e-13 PD=1.8e-06 PS=2.24496e-06 $X=6040 $Y=1185 $dt=0
M7 11 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=9e-14 AS=6.21542e-13 PD=9.7e-07 PS=3.8485e-06 $X=7495 $Y=660 $dt=0
M8 7 12 11 gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=2.26611e-13 AS=9e-14 PD=1.59158e-06 PS=9.7e-07 $X=8095 $Y=660 $dt=0
M9 10 13 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.32189e-13 PD=6.7e-07 PS=9.28421e-07 $X=8985 $Y=960 $dt=0
M10 gnd3i! 9 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.58966e-13 AS=5.25e-14 PD=1.9689e-06 PS=6.7e-07 $X=9585 $Y=960 $dt=0
M11 9 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.58966e-13 PD=1.8e-06 PS=1.9689e-06 $X=10355 $Y=1130 $dt=0
M12 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=7.60667e-13 PD=1.43e-06 PS=4.1722e-06 $X=11910 $Y=660 $dt=0
M13 gnd3i! 7 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=8.454e-13 AS=2.403e-13 PD=3.9e-06 PS=1.43e-06 $X=12800 $Y=660 $dt=0
M14 vdd3i! 8 16 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=6.82011e-13 AS=3.456e-13 PD=2.84211e-06 PS=2.4e-06 $X=620 $Y=2890 $dt=1
M15 20 16 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=7.35e-14 AS=3.97839e-13 PD=7.7e-07 PS=1.65789e-06 $X=1890 $Y=3400 $dt=1
M16 8 13 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.22795e-13 AS=7.35e-14 PD=9.06316e-07 PS=7.7e-07 $X=2540 $Y=3400 $dt=1
M17 19 12 8 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=1.375e-13 AS=3.21605e-13 PD=1.35e-06 PS=2.37368e-06 $X=3380 $Y=2720 $dt=1
M18 vdd3i! D 19 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=4.82459e-13 AS=1.375e-13 PD=2.50824e-06 PS=1.35e-06 $X=3930 $Y=2720 $dt=1
M19 13 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.78e-13 AS=3.15791e-13 PD=2.49e-06 PS=1.64176e-06 $X=4855 $Y=2720 $dt=1
M20 vdd3i! 13 12 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.24385e-13 AS=3.636e-13 PD=1.65561e-06 PS=2.45e-06 $X=6545 $Y=2670 $dt=1
M21 18 16 vdd3i! vdd3i! pe3i L=3e-07 W=1.15e-06 AD=1.4375e-13 AS=5.18115e-13 PD=1.4e-06 PS=2.64439e-06 $X=7495 $Y=2670 $dt=1
M22 7 13 18 vdd3i! pe3i L=3e-07 W=1.15e-06 AD=3.62506e-13 AS=1.4375e-13 PD=2.51975e-06 PS=1.4e-06 $X=8045 $Y=2670 $dt=1
M23 17 12 7 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.32394e-13 PD=6.7e-07 PS=9.20255e-07 $X=8915 $Y=3235 $dt=1
M24 vdd3i! 9 17 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=4.12999e-13 AS=5.25e-14 PD=1.6932e-06 PS=6.7e-07 $X=9465 $Y=3235 $dt=1
M25 9 7 vdd3i! vdd3i! pe3i L=3e-07 W=7.15e-07 AD=3.68225e-13 AS=7.03081e-13 PD=2.46e-06 PS=2.88248e-06 $X=10380 $Y=2410 $dt=1
M26 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.3865e-12 PD=1.95e-06 PS=5.68432e-06 $X=11960 $Y=2410 $dt=1
M27 vdd3i! 7 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.2851e-12 AS=3.807e-13 PD=5.04e-06 PS=1.95e-06 $X=12800 $Y=2410 $dt=1
.ends DFRQJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2JI3VX0 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 Q B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=7.244e-13 PD=9.6e-07 PS=4.14e-06 $X=500 $Y=1130 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=7.244e-13 AS=1.134e-13 PD=4.14e-06 PS=9.6e-07 $X=1390 $Y=1130 $dt=0
M2 7 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=9.298e-13 PD=1.1e-06 PS=4.68e-06 $X=720 $Y=2410 $dt=1
M3 Q A 7 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=1.0625e-13 PD=2.66e-06 PS=1.1e-06 $X=1270 $Y=2410 $dt=1
.ends NO2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN21JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.47e-13 PD=1.14e-06 PS=3.58e-06 $X=690 $Y=660 $dt=0
M1 Q A 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28413e-13 AS=1.1125e-13 PD=1.78572e-06 PS=1.14e-06 $X=1290 $Y=660 $dt=0
M2 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=6.369e-13 AS=2.45387e-13 PD=3.6e-06 PS=1.33428e-06 $X=2310 $Y=885 $dt=0
M3 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.371e-13 AS=6.768e-13 PD=2.03e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M4 9 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=4.371e-13 PD=1.95e-06 PS=2.03e-06 $X=1540 $Y=2410 $dt=1
M5 Q C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.614e-13 AS=3.807e-13 PD=3.9e-06 PS=1.95e-06 $X=2380 $Y=2410 $dt=1
.ends AN21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN22JI3VX1 vdd3i! gnd3i! B A Q C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 10 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.098e-13 PD=1.14e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 Q A 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=1260 $Y=660 $dt=0
M2 9 C Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.403e-13 PD=1.14e-06 PS=1.43e-06 $X=2150 $Y=660 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=8.082e-13 AS=1.1125e-13 PD=3.84e-06 PS=1.14e-06 $X=2750 $Y=660 $dt=0
M4 vdd3i! B 11 vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=4.29e-13 AS=6.0945e-13 PD=2.32213e-06 PS=3.77213e-06 $X=660 $Y=2410 $dt=1
M5 11 A vdd3i! vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=4.05825e-13 AS=4.29e-13 PD=2.06213e-06 PS=2.32213e-06 $X=1310 $Y=2410 $dt=1
M6 Q C 11 vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=2.9925e-13 AS=4.05825e-13 PD=1.92213e-06 PS=2.06213e-06 $X=2200 $Y=2410 $dt=1
M7 11 D Q vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=6.252e-13 AS=2.9925e-13 PD=3.77213e-06 PS=1.92213e-06 $X=3100 $Y=2410 $dt=1
.ends AN22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON211JI3VX1 vdd3i! gnd3i! B Q A C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 Q B 10 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.27987e-13 AS=4.20337e-13 PD=1.41536e-06 PS=2.75536e-06 $X=620 $Y=660 $dt=0
M1 10 A Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.30287e-13 AS=2.27987e-13 PD=1.43036e-06 PS=1.41536e-06 $X=1460 $Y=660 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=1.21188e-13 AS=2.30287e-13 PD=1.17536e-06 PS=1.43036e-06 $X=2350 $Y=660 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=4.20337e-13 AS=1.21188e-13 PD=2.75536e-06 PS=1.17536e-06 $X=2950 $Y=660 $dt=0
M4 11 B vdd3i! vdd3i! pe3i L=3e-07 W=1.38e-06 AD=1.725e-13 AS=9.388e-13 PD=1.63e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M5 Q A 11 vdd3i! pe3i L=3e-07 W=1.38e-06 AD=4.69617e-13 AS=1.725e-13 PD=2.38255e-06 PS=1.63e-06 $X=1245 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00049e-07 W=9.66924e-07 AD=4.25413e-13 AS=3.29046e-13 PD=2.34192e-06 PS=1.66938e-06 $X=2210 $Y=2410 $dt=1
M7 Q D vdd3i! vdd3i! pe3i L=3.00049e-07 W=9.66924e-07 AD=4.20162e-13 AS=4.25413e-13 PD=2.80192e-06 PS=2.34192e-06 $X=3000 $Y=2410 $dt=1
.ends ON211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EN2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EN2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=10 EP=5 FDC=10
M0 8 A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=620 $Y=980 $dt=0
M1 gnd3i! B 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=1220 $Y=980 $dt=0
M2 7 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=1.134e-13 PD=9.6e-07 PS=9.6e-07 $X=2110 $Y=980 $dt=0
M3 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.698e-13 AS=1.134e-13 PD=3.22e-06 PS=9.6e-07 $X=3000 $Y=980 $dt=0
M4 Q 9 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.058e-13 PD=1.8e-06 PS=1.82e-06 $X=4440 $Y=1020 $dt=0
M5 9 A vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=3.195e-13 AS=8.517e-13 PD=1.61e-06 PS=4.61e-06 $X=685 $Y=2410 $dt=1
M6 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=9e-07 AD=4.30855e-13 AS=3.195e-13 PD=1.83273e-06 PS=1.61e-06 $X=1695 $Y=2410 $dt=1
M7 10 A vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=6.22345e-13 PD=1.6e-06 PS=2.64727e-06 $X=2825 $Y=2520 $dt=1
M8 Q B 10 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=6.21324e-13 AS=1.95e-13 PD=2.52941e-06 PS=1.6e-06 $X=3425 $Y=2520 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=9.1e-07 AD=8.0675e-13 AS=4.34926e-13 PD=4.39e-06 PS=1.77059e-06 $X=4575 $Y=2520 $dt=1
.ends EN2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX0 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.892e-13 PD=8.1e-07 PS=3.54e-06 $X=670 $Y=990 $dt=0
M1 Q A 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.688e-13 AS=7e-14 PD=2.08e-06 PS=8.1e-07 $X=1270 $Y=990 $dt=0
M2 Q B vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=1.1114e-12 PD=1.24e-06 PS=4.94e-06 $X=550 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3e-07 W=7e-07 AD=1.1114e-12 AS=1.89e-13 PD=4.94e-06 PS=1.24e-06 $X=1390 $Y=2410 $dt=1
.ends NA2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX0                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX0 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=2
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=6.248e-13 PD=1.8e-06 PS=3.62e-06 $X=710 $Y=1130 $dt=0
M1 Q A vdd3i! vdd3i! pe3i L=3e-07 W=9.4e-07 AD=4.512e-13 AS=1.0092e-12 PD=2.84e-06 PS=4.76e-06 $X=760 $Y=2410 $dt=1
.ends INJI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRQJI3VX4                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRQJI3VX4 vdd3i! gnd3i! D C Q
*.DEVICECLIMB
** N=20 EP=5 FDC=32
M0 gnd3i! 9 16 gnd3i! ne3i L=3.5e-07 W=7.6e-07 AD=2.42427e-13 AS=3.648e-13 PD=1.67458e-06 PS=2.48e-06 $X=620 $Y=660 $dt=0
M1 15 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=6.09e-14 AS=1.33973e-13 PD=7.1e-07 PS=9.25424e-07 $X=1510 $Y=1000 $dt=0
M2 9 12 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.30725e-13 AS=6.09e-14 PD=9.3e-07 PS=7.1e-07 $X=2150 $Y=1000 $dt=0
M3 14 13 9 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=2.17875e-13 PD=9.5e-07 PS=1.55e-06 $X=3040 $Y=960 $dt=0
M4 gnd3i! D 14 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=6.04277e-13 AS=8.75e-14 PD=3.74159e-06 PS=9.5e-07 $X=3640 $Y=960 $dt=0
M5 gnd3i! C 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.62566e-13 AS=2.016e-13 PD=2.24496e-06 PS=1.8e-06 $X=5070 $Y=1295 $dt=0
M6 12 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.62566e-13 PD=1.8e-06 PS=2.24496e-06 $X=6040 $Y=1185 $dt=0
M7 11 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=9e-14 AS=6.21542e-13 PD=9.7e-07 PS=3.8485e-06 $X=7495 $Y=660 $dt=0
M8 8 12 11 gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=2.26611e-13 AS=9e-14 PD=1.59158e-06 PS=9.7e-07 $X=8095 $Y=660 $dt=0
M9 10 13 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.32189e-13 PD=6.7e-07 PS=9.28421e-07 $X=8985 $Y=960 $dt=0
M10 gnd3i! 7 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.98371e-13 AS=5.25e-14 PD=1.83685e-06 PS=6.7e-07 $X=9585 $Y=960 $dt=0
M11 7 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=3.29987e-13 AS=4.68868e-13 PD=2.26406e-06 PS=2.88647e-06 $X=10555 $Y=890 $dt=0
M12 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.32261e-13 PD=1.43e-06 PS=3.89237e-06 $X=12040 $Y=660 $dt=0
M13 gnd3i! 8 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=12930 $Y=660 $dt=0
M14 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=13820 $Y=660 $dt=0
M15 gnd3i! 8 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=14710 $Y=660 $dt=0
M16 vdd3i! 9 16 vdd3i! pe3i L=3e-07 W=1.11e-06 AD=9.09003e-13 AS=5.328e-13 PD=3.52588e-06 PS=3.18e-06 $X=620 $Y=2710 $dt=1
M17 20 16 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=7.35e-14 AS=3.43947e-13 PD=7.7e-07 PS=1.33412e-06 $X=1890 $Y=3400 $dt=1
M18 9 13 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.22795e-13 AS=7.35e-14 PD=9.06316e-07 PS=7.7e-07 $X=2540 $Y=3400 $dt=1
M19 19 12 9 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=1.375e-13 AS=3.21605e-13 PD=1.35e-06 PS=2.37368e-06 $X=3380 $Y=2720 $dt=1
M20 vdd3i! D 19 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=4.82459e-13 AS=1.375e-13 PD=2.50824e-06 PS=1.35e-06 $X=3930 $Y=2720 $dt=1
M21 13 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.78e-13 AS=3.15791e-13 PD=2.49e-06 PS=1.64176e-06 $X=4855 $Y=2720 $dt=1
M22 vdd3i! 13 12 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.24385e-13 AS=3.636e-13 PD=1.65561e-06 PS=2.45e-06 $X=6545 $Y=2670 $dt=1
M23 18 16 vdd3i! vdd3i! pe3i L=3e-07 W=1.15e-06 AD=1.4375e-13 AS=5.18115e-13 PD=1.4e-06 PS=2.64439e-06 $X=7495 $Y=2670 $dt=1
M24 8 13 18 vdd3i! pe3i L=3e-07 W=1.15e-06 AD=3.62506e-13 AS=1.4375e-13 PD=2.51975e-06 PS=1.4e-06 $X=8045 $Y=2670 $dt=1
M25 17 12 8 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.32394e-13 PD=6.7e-07 PS=9.20255e-07 $X=8915 $Y=3235 $dt=1
M26 vdd3i! 7 17 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=2.19743e-13 AS=5.25e-14 PD=1.10393e-06 PS=6.7e-07 $X=9465 $Y=3235 $dt=1
M27 7 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.2615e-13 AS=7.37707e-13 PD=3.85e-06 PS=3.70607e-06 $X=10410 $Y=2410 $dt=1
M28 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.2586e-12 PD=1.95e-06 PS=4.99e-06 $X=12240 $Y=2410 $dt=1
M29 vdd3i! 8 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=3.807e-13 PD=1.95e-06 PS=1.95e-06 $X=13080 $Y=2410 $dt=1
M30 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=3.807e-13 PD=1.95e-06 PS=1.95e-06 $X=13920 $Y=2410 $dt=1
M31 vdd3i! 8 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=3.807e-13 PD=3.78e-06 PS=1.95e-06 $X=14760 $Y=2410 $dt=1
.ends DFRQJI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRQJI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRQJI3VX1 vdd3i! gnd3i! D C Q
*.DEVICECLIMB
** N=20 EP=5 FDC=26
M0 gnd3i! 8 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=2.016e-13 PD=9.6e-07 PS=1.8e-06 $X=620 $Y=1000 $dt=0
M1 15 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=6.09e-14 AS=1.134e-13 PD=7.1e-07 PS=9.6e-07 $X=1510 $Y=1000 $dt=0
M2 8 12 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.30725e-13 AS=6.09e-14 PD=9.3e-07 PS=7.1e-07 $X=2150 $Y=1000 $dt=0
M3 14 13 8 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=2.17875e-13 PD=9.5e-07 PS=1.55e-06 $X=3040 $Y=960 $dt=0
M4 gnd3i! D 14 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=6.04277e-13 AS=8.75e-14 PD=3.74159e-06 PS=9.5e-07 $X=3640 $Y=960 $dt=0
M5 gnd3i! C 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.62566e-13 AS=2.016e-13 PD=2.24496e-06 PS=1.8e-06 $X=5070 $Y=1295 $dt=0
M6 12 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.62566e-13 PD=1.8e-06 PS=2.24496e-06 $X=6040 $Y=1185 $dt=0
M7 11 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=9e-14 AS=6.21542e-13 PD=9.7e-07 PS=3.8485e-06 $X=7495 $Y=660 $dt=0
M8 7 12 11 gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=2.26611e-13 AS=9e-14 PD=1.59158e-06 PS=9.7e-07 $X=8095 $Y=660 $dt=0
M9 10 13 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.32189e-13 PD=6.7e-07 PS=9.28421e-07 $X=8985 $Y=960 $dt=0
M10 gnd3i! 9 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.58966e-13 AS=5.25e-14 PD=1.9689e-06 PS=6.7e-07 $X=9585 $Y=960 $dt=0
M11 9 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.58966e-13 PD=1.8e-06 PS=1.9689e-06 $X=10355 $Y=1130 $dt=0
M12 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=7.60667e-13 PD=2.74e-06 PS=4.1722e-06 $X=11910 $Y=660 $dt=0
M13 vdd3i! 8 16 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=6.82011e-13 AS=3.456e-13 PD=2.84211e-06 PS=2.4e-06 $X=620 $Y=2890 $dt=1
M14 20 16 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=7.35e-14 AS=3.97839e-13 PD=7.7e-07 PS=1.65789e-06 $X=1890 $Y=3400 $dt=1
M15 8 13 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.22795e-13 AS=7.35e-14 PD=9.06316e-07 PS=7.7e-07 $X=2540 $Y=3400 $dt=1
M16 19 12 8 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=1.375e-13 AS=3.21605e-13 PD=1.35e-06 PS=2.37368e-06 $X=3380 $Y=2720 $dt=1
M17 vdd3i! D 19 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=4.82459e-13 AS=1.375e-13 PD=2.50824e-06 PS=1.35e-06 $X=3930 $Y=2720 $dt=1
M18 13 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.78e-13 AS=3.15791e-13 PD=2.49e-06 PS=1.64176e-06 $X=4855 $Y=2720 $dt=1
M19 vdd3i! 13 12 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.24385e-13 AS=3.636e-13 PD=1.65561e-06 PS=2.45e-06 $X=6545 $Y=2670 $dt=1
M20 18 16 vdd3i! vdd3i! pe3i L=3e-07 W=1.15e-06 AD=1.4375e-13 AS=5.18115e-13 PD=1.4e-06 PS=2.64439e-06 $X=7495 $Y=2670 $dt=1
M21 7 13 18 vdd3i! pe3i L=3e-07 W=1.15e-06 AD=3.62506e-13 AS=1.4375e-13 PD=2.51975e-06 PS=1.4e-06 $X=8045 $Y=2670 $dt=1
M22 17 12 7 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.32394e-13 PD=6.7e-07 PS=9.20255e-07 $X=8915 $Y=3235 $dt=1
M23 vdd3i! 9 17 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=4.12999e-13 AS=5.25e-14 PD=1.6932e-06 PS=6.7e-07 $X=9465 $Y=3235 $dt=1
M24 9 7 vdd3i! vdd3i! pe3i L=3e-07 W=7.15e-07 AD=3.68225e-13 AS=7.03081e-13 PD=2.46e-06 PS=2.88248e-06 $X=10380 $Y=2410 $dt=1
M25 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.3865e-12 PD=3.78e-06 PS=5.68432e-06 $X=11960 $Y=2410 $dt=1
.ends DFRQJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP25JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP25JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=12
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=3990 $Y=660 $dt=0
M3 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=6470 $Y=660 $dt=0
M4 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=8950 $Y=660 $dt=0
M5 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=4.312e-13 AS=2.376e-13 PD=2.74e-06 PS=1.42e-06 $X=11430 $Y=660 $dt=0
M6 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=6.312e-13 PD=1.855e-06 PS=3.59e-06 $X=620 $Y=2505 $dt=1
M7 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=3090 $Y=2505 $dt=1
M8 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=5560 $Y=2505 $dt=1
M9 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=8030 $Y=2505 $dt=1
M10 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.84638e-13 AS=3.5505e-13 PD=1.9e-06 PS=1.855e-06 $X=10500 $Y=2505 $dt=1
M11 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.84638e-13 PD=3.91e-06 PS=1.9e-06 $X=13015 $Y=2505 $dt=1
.ends DECAP25JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP10JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP10JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=6
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.445e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.445e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=3495 $Y=660 $dt=0
M3 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.425e-06 W=1.315e-06 AD=3.5505e-13 AS=8.308e-13 PD=1.855e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M4 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.425e-06 W=1.315e-06 AD=3.71488e-13 AS=3.5505e-13 PD=1.88e-06 PS=1.855e-06 $X=2625 $Y=2505 $dt=1
M5 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.71488e-13 PD=3.91e-06 PS=1.88e-06 $X=4615 $Y=2505 $dt=1
.ends DECAP10JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP7JI3V                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP7JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=4
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.75e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.71e-06 W=1.315e-06 AD=3.87925e-13 AS=8.308e-13 PD=1.905e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M3 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.237e-13 AS=3.87925e-13 PD=3.86e-06 PS=1.905e-06 $X=2960 $Y=2505 $dt=1
.ends DECAP7JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP15JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP15JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=8
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.42e-13 AS=4.224e-13 PD=1.43e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=2.42e-13 AS=2.42e-13 PD=1.43e-06 PS=1.43e-06 $X=1520 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=2.376e-13 AS=2.42e-13 PD=1.42e-06 PS=1.43e-06 $X=3780 $Y=660 $dt=0
M3 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=6030 $Y=660 $dt=0
M4 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.5505e-13 AS=8.308e-13 PD=1.855e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M5 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=2900 $Y=2505 $dt=1
M6 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.78063e-13 AS=3.5505e-13 PD=1.89e-06 PS=1.855e-06 $X=5140 $Y=2505 $dt=1
M7 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.78063e-13 PD=3.91e-06 PS=1.89e-06 $X=7415 $Y=2505 $dt=1
.ends DECAP15JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP5JI3V                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP5JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=2
M0 gnd3i! 5 4 gnd3i! ne3i L=1.48e-06 W=8.3e-07 AD=5.786e-13 AS=4.568e-13 PD=3.4e-06 PS=2.82e-06 $X=660 $Y=660 $dt=0
M1 5 4 vdd3i! vdd3i! pe3i L=1.46e-06 W=1.36e-06 AD=7.564e-13 AS=8.542e-13 PD=3.9e-06 PS=4.46e-06 $X=660 $Y=2460 $dt=1
.ends DECAP5JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: counter                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt counter 1 2 3 out<7> out<6> enable out<2> out<3> out<5> out<4>
+ reset out<1> out<0> clk
** N=62 EP=14 FDC=711
X287 2 3 55 18 BUJI3VX2 $T=24080 32480 1 0 $X=23650 $Y=27360
X288 2 3 30 out<0> BUJI3VX2 $T=50960 14560 1 0 $X=50530 $Y=9440
X289 2 3 15 16 BUJI3VX0 $T=15120 50400 1 0 $X=14690 $Y=45280
X290 2 3 41 34 BUJI3VX16 $T=11200 50400 0 0 $X=10770 $Y=49760
X291 2 3 42 46 DLY1JI3VX1 $T=18480 14560 0 0 $X=18050 $Y=13920
X292 2 3 44 43 DLY1JI3VX1 $T=51520 41440 1 0 $X=51090 $Y=36320
X293 2 3 enable 19 DLY2JI3VX1 $T=27440 50400 0 0 $X=27010 $Y=49760
X294 2 3 reset 20 DLY2JI3VX1 $T=39200 50400 0 0 $X=38770 $Y=49760
X295 2 3 23 36 DLY2JI3VX1 $T=49280 32480 0 0 $X=48850 $Y=31840
X296 2 3 51 39 DLY2JI3VX1 $T=49840 32480 1 0 $X=49410 $Y=27360
X297 2 3 54 31 DLY2JI3VX1 $T=53200 14560 0 0 $X=52770 $Y=13920
X298 2 3 40 17 BUJI3VX1 $T=20160 41440 0 0 $X=19730 $Y=40800
X299 2 3 clk 40 BUJI3VX1 $T=56000 50400 0 0 $X=55570 $Y=49760
X300 2 3 18 17 out<7> DFRQJI3VX2 $T=31360 23520 1 180 $X=16930 $Y=22880
X301 2 3 16 17 out<6> DFRQJI3VX2 $T=17920 50400 1 0 $X=17490 $Y=45280
X302 2 3 46 17 out<3> DFRQJI3VX2 $T=18480 23520 1 0 $X=18050 $Y=18400
X303 2 3 36 17 out<2> DFRQJI3VX2 $T=45920 23520 1 180 $X=31490 $Y=22880
X304 2 3 34 17 out<5> DFRQJI3VX2 $T=34720 50400 1 0 $X=34290 $Y=45280
X305 2 3 43 17 out<4> DFRQJI3VX2 $T=37520 41440 1 0 $X=37090 $Y=36320
X306 2 3 47 55 20 NO2JI3VX0 $T=29680 32480 0 180 $X=27010 $Y=27360
X307 2 3 56 51 20 NO2JI3VX0 $T=49840 32480 0 180 $X=47170 $Y=27360
X308 2 3 57 33 15 20 AN21JI3VX1 $T=26880 41440 1 180 $X=23090 $Y=40800
X309 2 3 58 21 42 20 AN21JI3VX1 $T=27440 14560 1 180 $X=23650 $Y=13920
X310 2 3 59 53 23 20 AN21JI3VX1 $T=41440 23520 0 180 $X=37650 $Y=18400
X311 2 3 27 37 41 20 AN21JI3VX1 $T=40320 41440 0 0 $X=39890 $Y=40800
X312 2 3 28 52 44 20 AN21JI3VX1 $T=42560 32480 0 0 $X=42130 $Y=31840
X313 2 3 60 38 54 20 AN21JI3VX1 $T=45920 14560 0 0 $X=45490 $Y=13920
X314 2 3 19 61 47 out<7> 25 AN22JI3VX1 $T=27440 32480 0 0 $X=27010 $Y=31840
X315 2 3 out<6> 33 62 32 19 ON211JI3VX1 $T=29120 41440 0 180 $X=24770 $Y=36320
X316 2 3 out<3> 21 49 35 19 ON211JI3VX1 $T=35280 14560 1 180 $X=30930 $Y=13920
X317 2 3 out<5> 37 22 50 19 ON211JI3VX1 $T=31360 41440 0 0 $X=30930 $Y=40800
X318 2 3 out<2> 53 26 24 19 ON211JI3VX1 $T=38640 14560 1 0 $X=38210 $Y=9440
X319 2 3 out<4> 52 48 45 19 ON211JI3VX1 $T=38640 32480 0 0 $X=38210 $Y=31840
X320 2 3 out<1> 38 out<0> 29 19 ON211JI3VX1 $T=43680 14560 1 0 $X=43250 $Y=9440
X321 2 3 out<7> 32 61 EN2JI3VX0 $T=20720 32480 0 0 $X=20290 $Y=31840
X322 2 3 19 30 56 EN2JI3VX0 $T=42000 32480 1 0 $X=41570 $Y=27360
X323 2 3 out<6> 32 62 NA2JI3VX0 $T=21840 41440 1 0 $X=21410 $Y=36320
X324 2 3 25 57 out<6> NA2JI3VX0 $T=30240 41440 1 180 $X=27570 $Y=40800
X325 2 3 25 58 out<3> NA2JI3VX0 $T=28560 14560 0 0 $X=28130 $Y=13920
X326 2 3 out<3> 35 49 NA2JI3VX0 $T=29680 14560 1 0 $X=29250 $Y=9440
X327 2 3 out<4> 45 48 NA2JI3VX0 $T=34720 32480 0 180 $X=32050 $Y=27360
X328 2 3 out<5> 50 22 NA2JI3VX0 $T=34720 41440 0 180 $X=32050 $Y=36320
X329 2 3 out<2> 24 26 NA2JI3VX0 $T=39200 14560 0 0 $X=38770 $Y=13920
X330 2 3 25 59 out<2> NA2JI3VX0 $T=41440 23520 1 0 $X=41010 $Y=18400
X331 2 3 25 60 out<1> NA2JI3VX0 $T=42560 14560 0 0 $X=42130 $Y=13920
X332 2 3 25 27 out<5> NA2JI3VX0 $T=45920 41440 1 180 $X=43250 $Y=40800
X333 2 3 25 28 out<4> NA2JI3VX0 $T=49280 32480 1 180 $X=46610 $Y=31840
X334 2 3 out<1> 29 30 NA2JI3VX0 $T=50960 14560 0 0 $X=50530 $Y=13920
X335 2 3 50 62 INJI3VX0 $T=31920 41440 0 180 $X=29810 $Y=36320
X336 2 3 24 49 INJI3VX0 $T=34720 14560 0 180 $X=32610 $Y=9440
X337 2 3 35 48 INJI3VX0 $T=35280 23520 0 180 $X=33170 $Y=18400
X338 2 3 45 22 INJI3VX0 $T=35280 32480 1 180 $X=33170 $Y=31840
X339 2 3 19 25 INJI3VX0 $T=47600 41440 1 180 $X=45490 $Y=40800
X340 2 3 29 26 INJI3VX0 $T=49280 14560 0 180 $X=47170 $Y=9440
X341 2 3 31 17 out<1> DFRQJI3VX4 $T=44240 23520 1 0 $X=43810 $Y=18400
X342 2 3 39 17 30 DFRQJI3VX1 $T=45920 23520 0 0 $X=45490 $Y=22880
X343 2 3 DECAP25JI3V $T=10080 14560 1 0 $X=9650 $Y=9440
X344 2 3 DECAP10JI3V $T=10080 23520 0 0 $X=9650 $Y=22880
X345 2 3 DECAP10JI3V $T=10080 41440 0 0 $X=9650 $Y=40800
X346 2 3 DECAP10JI3V $T=24080 14560 1 0 $X=23650 $Y=9440
X347 2 3 DECAP10JI3V $T=52080 50400 1 180 $X=46050 $Y=49760
X348 2 3 DECAP10JI3V $T=54320 14560 1 0 $X=53890 $Y=9440
X349 2 3 DECAP7JI3V $T=10080 32480 0 0 $X=9650 $Y=31840
X350 2 3 DECAP7JI3V $T=10080 41440 1 0 $X=9650 $Y=36320
X351 2 3 DECAP7JI3V $T=10080 50400 1 0 $X=9650 $Y=45280
X352 2 3 DECAP7JI3V $T=14000 32480 0 0 $X=13570 $Y=31840
X353 2 3 DECAP7JI3V $T=14000 41440 1 0 $X=13570 $Y=36320
X354 2 3 DECAP7JI3V $T=17920 41440 1 0 $X=17490 $Y=36320
X355 2 3 DECAP7JI3V $T=34720 14560 1 0 $X=34290 $Y=9440
X356 2 3 DECAP7JI3V $T=47600 41440 0 0 $X=47170 $Y=40800
X357 2 3 DECAP7JI3V $T=48720 50400 1 0 $X=48290 $Y=45280
X358 2 3 DECAP7JI3V $T=51520 41440 0 0 $X=51090 $Y=40800
X359 2 3 DECAP7JI3V $T=52080 50400 0 0 $X=51650 $Y=49760
X360 2 3 DECAP7JI3V $T=52640 50400 1 0 $X=52210 $Y=45280
X361 2 3 DECAP7JI3V $T=55440 41440 0 0 $X=55010 $Y=40800
X362 2 3 DECAP7JI3V $T=56560 32480 0 0 $X=56130 $Y=31840
X363 2 3 DECAP7JI3V $T=56560 50400 1 0 $X=56130 $Y=45280
X364 2 3 DECAP7JI3V $T=57120 32480 1 0 $X=56690 $Y=27360
X365 2 3 DECAP7JI3V $T=57120 41440 1 0 $X=56690 $Y=36320
X366 2 3 DECAP7JI3V $T=59360 41440 0 0 $X=58930 $Y=40800
X367 2 3 DECAP15JI3V $T=10080 14560 0 0 $X=9650 $Y=13920
X368 2 3 DECAP15JI3V $T=10080 23520 1 0 $X=9650 $Y=18400
X369 2 3 DECAP15JI3V $T=10080 32480 1 0 $X=9650 $Y=27360
X370 2 3 DECAP5JI3V $T=15680 41440 0 0 $X=15250 $Y=40800
X371 2 3 DECAP5JI3V $T=18480 32480 1 0 $X=18050 $Y=27360
X372 2 3 DECAP5JI3V $T=31920 50400 1 0 $X=31490 $Y=45280
X373 2 3 DECAP5JI3V $T=34720 41440 1 0 $X=34290 $Y=36320
X374 2 3 DECAP5JI3V $T=34720 50400 0 0 $X=34290 $Y=49760
X375 2 3 DECAP5JI3V $T=35280 23520 1 0 $X=34850 $Y=18400
X376 2 3 DECAP5JI3V $T=58800 23520 0 0 $X=58370 $Y=22880
X377 2 3 DECAP5JI3V $T=58800 50400 0 0 $X=58370 $Y=49760
X378 2 3 DECAP5JI3V $T=60480 14560 0 0 $X=60050 $Y=13920
X379 2 3 DECAP5JI3V $T=60480 32480 0 0 $X=60050 $Y=31840
X380 2 3 DECAP5JI3V $T=60480 50400 1 0 $X=60050 $Y=45280
D0 1 2 p_ddnwmv AREA=4.92445e-09 PJ=0.0002812 perimeter=0.0002812 $X=-570 $Y=-570 $dt=2
D1 3 2 p_dipdnwmv AREA=2.16064e-10 PJ=0.000116905 perimeter=0.000116905 $X=9650 $Y=12580 $dt=3
D2 3 2 p_dipdnwmv AREA=2.19665e-10 PJ=0.000117426 perimeter=0.000117426 $X=20170 $Y=48160 $dt=3
D3 3 2 p_dipdnwmv AREA=2.22073e-10 PJ=0.000117878 perimeter=0.000117878 $X=20730 $Y=21280 $dt=3
D4 3 2 p_dipdnwmv AREA=2.16467e-10 PJ=0.000116691 perimeter=0.000116691 $X=50340 $Y=30270 $dt=3
D5 3 2 p_dipdnwmv AREA=2.16468e-10 PJ=0.000116948 perimeter=0.000116948 $X=51970 $Y=39190 $dt=3
.ends counter

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: counter_lvs                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt counter_lvs gndd vddd vsub
** N=14 EP=3 FDC=711
X0 vsub vddd gndd 4 5 6 7 8 9 10
+ 11 12 13 14 counter $T=4235 4350 0 0 $X=2795 $Y=2910
.ends counter_lvs
