
wire \gnd3i! ;

wire \vdd3i! ;

wire \gnd! ;
