* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ioring3                                      *
* Netlisted  : Sat Feb 10 19:20:57 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3i) nemi ndiff(D) p1trm(G) ndiff(S) pwitrm(B)
*.DEVTMPLT 1 MP(pe3i) pemi pdiff(D) p1trm(G) pdiff(S) dnwtrm(B)
*.DEVTMPLT 2 D(ddnwmv) d_ddnwmv bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 3 D(p_ddnwmv) p_ddnwmv bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 4 D(dipdnwmv) d_dipwmv pwitrm(POS) dnwtrm(NEG)
*.DEVTMPLT 5 R(rdn3) rdnm_gi ndiff(POS) ndiff(NEG) pwitrm(SUB)
*.DEVTMPLT 6 R(rdp3) rdpm pdiff(POS) pdiff(NEG) nwtrm(SUB)
*.DEVTMPLT 7 R(rdp3) rdpmi pdiff(POS) pdiff(NEG) dnwtrm(SUB)
*.DEVTMPLT 8 R(rdp3) rdpm_gi pdiff(POS) pdiff(NEG) dnwtrm(SUB)
*.DEVTMPLT 9 D(dn3) d_dnmi1 pwitrm(POS) ndiff(NEG)
*.DEVTMPLT 10 D(dp3) d_dpm pdiff(POS) nwtrm(NEG)
*.DEVTMPLT 11 D(p_dp3) p_dpm pdiff(POS) nwtrm(NEG)
*.DEVTMPLT 12 D(p_dp3) p_dpmi1 pdiff(POS) dnwtrm(NEG)
*.DEVTMPLT 13 D(p_dnw3) p_dnwm bulk(POS) nwtrm(NEG)
*.DEVTMPLT 14 R(rpp1) rpp1_2 p1trm(POS) p1trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_pe3isb_pc                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_pe3isb_pc 2 3 6 7
*.DEVICECLIMB
** N=10 EP=4 FDC=3
R0 7 3 L=2.15e-06 W=3e-05 $[rdp3] $SUB=2 $X=1000 $Y=1825 $dt=8
R1 3 6 L=2.15e-06 W=3e-05 $[rdp3] $SUB=2 $X=3805 $Y=1825 $dt=8
D2 3 2 p_dp3 AREA=1.98e-11 PJ=1.32e-06 perimeter=1.32e-06 $X=3145 $Y=1825 $dt=12
.ends jio_pe3isb_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_ne3isbg_pc                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_ne3isbg_pc 2 3 5 6
*.DEVICECLIMB
** N=9 EP=4 FDC=3
R0 5 3 L=3.35e-06 W=3e-05 $[rdn3] $SUB=2 $X=955 $Y=1825 $dt=5
R1 3 6 L=3.35e-06 W=3e-05 $[rdn3] $SUB=2 $X=4960 $Y=1825 $dt=5
D2 2 3 dn3 AREA=1.98e-11 PJ=1.32e-06 perimeter=1.32e-06 $X=4300 $Y=1825 $dt=9
.ends jio_ne3isbg_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: PSUBPADPC                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt PSUBPADPC PSUB GNDOI VDDOI VDD3I GNDI VDDRI GNDRI
** N=65 EP=7 FDC=149
X1174 VDDOI PSUB 37 36 jio_pe3isb_pc $T=14365 150990 1 180 $X=6700 $Y=149060
X1175 VDDOI PSUB 35 34 jio_pe3isb_pc $T=14365 184790 1 180 $X=6700 $Y=182860
X1176 VDDOI PSUB 45 44 jio_pe3isb_pc $T=20965 150990 1 180 $X=13300 $Y=149060
X1177 VDDOI PSUB 43 42 jio_pe3isb_pc $T=20965 184790 1 180 $X=13300 $Y=182860
X1178 VDDOI PSUB 41 40 jio_pe3isb_pc $T=27565 150990 1 180 $X=19900 $Y=149060
X1179 VDDOI PSUB 39 38 jio_pe3isb_pc $T=27565 184790 1 180 $X=19900 $Y=182860
X1180 VDDOI PSUB 49 48 jio_pe3isb_pc $T=34165 150990 1 180 $X=26500 $Y=149060
X1181 VDDOI PSUB 47 46 jio_pe3isb_pc $T=34165 184790 1 180 $X=26500 $Y=182860
X1182 VDDOI PSUB 57 56 jio_pe3isb_pc $T=35835 150990 0 0 $X=35120 $Y=149060
X1183 VDDOI PSUB 55 54 jio_pe3isb_pc $T=35835 184790 0 0 $X=35120 $Y=182860
X1184 VDDOI PSUB 53 52 jio_pe3isb_pc $T=42435 150990 0 0 $X=41720 $Y=149060
X1185 VDDOI PSUB 51 50 jio_pe3isb_pc $T=42435 184790 0 0 $X=41720 $Y=182860
X1186 VDDOI PSUB 65 64 jio_pe3isb_pc $T=49035 150990 0 0 $X=48320 $Y=149060
X1187 VDDOI PSUB 63 62 jio_pe3isb_pc $T=49035 184790 0 0 $X=48320 $Y=182860
X1188 VDDOI PSUB 61 60 jio_pe3isb_pc $T=55635 150990 0 0 $X=54920 $Y=149060
X1189 VDDOI PSUB 59 58 jio_pe3isb_pc $T=55635 184790 0 0 $X=54920 $Y=182860
X1458 PSUB GNDOI 12 13 jio_ne3isbg_pc $T=16420 75080 1 180 $X=6100 $Y=74005
X1459 PSUB GNDOI 10 11 jio_ne3isbg_pc $T=16420 108880 1 180 $X=6100 $Y=107805
X1460 PSUB GNDOI 16 17 jio_ne3isbg_pc $T=25420 75080 1 180 $X=15100 $Y=74005
X1461 PSUB GNDOI 14 15 jio_ne3isbg_pc $T=25420 108880 1 180 $X=15100 $Y=107805
X1462 PSUB GNDOI 24 25 jio_ne3isbg_pc $T=34420 75080 1 180 $X=24100 $Y=74005
X1463 PSUB GNDOI 22 23 jio_ne3isbg_pc $T=34420 108880 1 180 $X=24100 $Y=107805
X1464 PSUB GNDOI 20 21 jio_ne3isbg_pc $T=35580 75080 0 0 $X=34520 $Y=74005
X1465 PSUB GNDOI 18 19 jio_ne3isbg_pc $T=35580 108880 0 0 $X=34520 $Y=107805
X1466 PSUB GNDOI 28 29 jio_ne3isbg_pc $T=44580 75080 0 0 $X=43520 $Y=74005
X1467 PSUB GNDOI 26 27 jio_ne3isbg_pc $T=44580 108880 0 0 $X=43520 $Y=107805
X1468 PSUB GNDOI 32 33 jio_ne3isbg_pc $T=53580 75080 0 0 $X=52520 $Y=74005
X1469 PSUB GNDOI 30 31 jio_ne3isbg_pc $T=53580 108880 0 0 $X=52520 $Y=107805
M0 13 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.89e-11 PD=6.001e-05 PS=6.126e-05 $X=7710 $Y=76905 $dt=0
M1 11 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.89e-11 PD=6.001e-05 PS=6.126e-05 $X=7710 $Y=110705 $dt=0
M2 PSUB 9 12 PSUB ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=15470 $Y=76905 $dt=0
M3 PSUB 9 10 PSUB ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=15470 $Y=110705 $dt=0
M4 17 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=16710 $Y=76905 $dt=0
M5 15 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=16710 $Y=110705 $dt=0
M6 PSUB 9 16 PSUB ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=24470 $Y=76905 $dt=0
M7 PSUB 9 14 PSUB ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=24470 $Y=110705 $dt=0
M8 25 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=25710 $Y=76905 $dt=0
M9 23 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=25710 $Y=110705 $dt=0
M10 PSUB 9 24 PSUB ne3i L=4e-07 W=3e-05 AD=3.39e-11 AS=1.5e-13 PD=3.226e-05 PS=6.001e-05 $X=33470 $Y=76905 $dt=0
M11 PSUB 9 22 PSUB ne3i L=4e-07 W=3e-05 AD=3.39e-11 AS=1.5e-13 PD=3.226e-05 PS=6.001e-05 $X=33470 $Y=110705 $dt=0
M12 20 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=3.39e-11 PD=6.001e-05 PS=3.226e-05 $X=36130 $Y=76905 $dt=0
M13 18 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=3.39e-11 PD=6.001e-05 PS=3.226e-05 $X=36130 $Y=110705 $dt=0
M14 PSUB 9 21 PSUB ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=43890 $Y=76905 $dt=0
M15 PSUB 9 19 PSUB ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=43890 $Y=110705 $dt=0
M16 28 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=45130 $Y=76905 $dt=0
M17 26 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=45130 $Y=110705 $dt=0
M18 PSUB 9 29 PSUB ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=52890 $Y=76905 $dt=0
M19 PSUB 9 27 PSUB ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=52890 $Y=110705 $dt=0
M20 32 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=54130 $Y=76905 $dt=0
M21 30 9 PSUB PSUB ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=54130 $Y=110705 $dt=0
M22 PSUB 9 33 PSUB ne3i L=4e-07 W=3e-05 AD=1.89e-11 AS=1.5e-13 PD=6.126e-05 PS=6.001e-05 $X=61890 $Y=76905 $dt=0
M23 PSUB 9 31 PSUB ne3i L=4e-07 W=3e-05 AD=1.89e-11 AS=1.5e-13 PD=6.126e-05 PS=6.001e-05 $X=61890 $Y=110705 $dt=0
M24 37 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=8060 $Y=152815 $dt=1
M25 35 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=8060 $Y=186615 $dt=1
M26 VDDOI 8 36 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=13370 $Y=152815 $dt=1
M27 VDDOI 8 34 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=13370 $Y=186615 $dt=1
M28 45 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=14660 $Y=152815 $dt=1
M29 43 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=14660 $Y=186615 $dt=1
M30 VDDOI 8 44 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=19970 $Y=152815 $dt=1
M31 VDDOI 8 42 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=19970 $Y=186615 $dt=1
M32 41 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=21260 $Y=152815 $dt=1
M33 39 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=21260 $Y=186615 $dt=1
M34 VDDOI 8 40 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=26570 $Y=152815 $dt=1
M35 VDDOI 8 38 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=26570 $Y=186615 $dt=1
M36 49 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=27860 $Y=152815 $dt=1
M37 47 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=27860 $Y=186615 $dt=1
M38 VDDOI 8 48 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=33170 $Y=152815 $dt=1
M39 VDDOI 8 46 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=33170 $Y=186615 $dt=1
M40 56 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=36480 $Y=152815 $dt=1
M41 54 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=36480 $Y=186615 $dt=1
M42 VDDOI 8 57 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=41790 $Y=152815 $dt=1
M43 VDDOI 8 55 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=41790 $Y=186615 $dt=1
M44 52 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=43080 $Y=152815 $dt=1
M45 50 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=43080 $Y=186615 $dt=1
M46 VDDOI 8 53 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=48390 $Y=152815 $dt=1
M47 VDDOI 8 51 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=48390 $Y=186615 $dt=1
M48 64 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=49680 $Y=152815 $dt=1
M49 62 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=49680 $Y=186615 $dt=1
M50 VDDOI 8 65 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=54990 $Y=152815 $dt=1
M51 VDDOI 8 63 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=54990 $Y=186615 $dt=1
M52 60 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=56280 $Y=152815 $dt=1
M53 58 8 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=56280 $Y=186615 $dt=1
M54 VDDOI 8 61 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=61590 $Y=152815 $dt=1
M55 VDDOI 8 59 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=61590 $Y=186615 $dt=1
D56 PSUB GNDOI ddnwmv AREA=4.69976e-09 PJ=0.00027464 perimeter=0.00027464 $X=2570 $Y=72575 $dt=2
D57 PSUB VDDOI p_ddnwmv AREA=4.5084e-09 PJ=0.00026872 perimeter=0.00026872 $X=2500 $Y=150035 $dt=3
D58 PSUB GNDOI dipdnwmv AREA=4.16648e-09 PJ=0.00025864 perimeter=0.00025864 $X=4570 $Y=74575 $dt=4
R59 8 VDDOI L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=VDDOI $X=4475 $Y=153720 $dt=7
R60 9 PSUB L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=VDDOI $X=65085 $Y=153720 $dt=7
D61 8 VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=4475 $Y=152700 $dt=12
D62 VDDOI VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=4475 $Y=157020 $dt=12
D63 9 VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=65085 $Y=152700 $dt=12
D64 PSUB VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=65085 $Y=157020 $dt=12
.ends PSUBPADPC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_ne3isb_pc                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_ne3isb_pc 2 3 6 7
*.DEVICECLIMB
** N=10 EP=4 FDC=3
R0 6 3 L=3.35e-06 W=3e-05 $[rdn3] $SUB=2 $X=955 $Y=1825 $dt=5
R1 3 7 L=3.35e-06 W=3e-05 $[rdn3] $SUB=2 $X=4960 $Y=1825 $dt=5
D2 2 3 dn3 AREA=1.98e-11 PJ=1.32e-06 perimeter=1.32e-06 $X=4300 $Y=1825 $dt=9
.ends jio_ne3isb_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_base_ntrc_pc                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_base_ntrc_pc 1 2 3 4 5
** N=29 EP=5 FDC=62
X100 2 4 8 9 jio_ne3isb_pc $T=16420 75080 1 180 $X=6100 $Y=73130
X101 2 4 6 7 jio_ne3isb_pc $T=16420 108880 1 180 $X=6100 $Y=106930
X102 2 4 12 13 jio_ne3isb_pc $T=25420 75080 1 180 $X=15100 $Y=73130
X103 2 4 10 11 jio_ne3isb_pc $T=25420 108880 1 180 $X=15100 $Y=106930
X104 2 4 16 17 jio_ne3isb_pc $T=34420 75080 1 180 $X=24100 $Y=73130
X105 2 4 14 15 jio_ne3isb_pc $T=34420 108880 1 180 $X=24100 $Y=106930
X106 2 4 20 21 jio_ne3isb_pc $T=35580 75080 0 0 $X=34520 $Y=73130
X107 2 4 18 19 jio_ne3isb_pc $T=35580 108880 0 0 $X=34520 $Y=106930
X108 2 4 24 25 jio_ne3isb_pc $T=44580 75080 0 0 $X=43520 $Y=73130
X109 2 4 22 23 jio_ne3isb_pc $T=44580 108880 0 0 $X=43520 $Y=106930
X110 2 4 28 29 jio_ne3isb_pc $T=53580 75080 0 0 $X=52520 $Y=73130
X111 2 4 26 27 jio_ne3isb_pc $T=53580 108880 0 0 $X=52520 $Y=106930
M0 9 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.89e-11 PD=6.001e-05 PS=6.126e-05 $X=7710 $Y=76905 $dt=0
M1 7 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.89e-11 PD=6.001e-05 PS=6.126e-05 $X=7710 $Y=110705 $dt=0
M2 2 3 8 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=15470 $Y=76905 $dt=0
M3 2 3 6 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=15470 $Y=110705 $dt=0
M4 13 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=16710 $Y=76905 $dt=0
M5 11 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=16710 $Y=110705 $dt=0
M6 2 3 12 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=24470 $Y=76905 $dt=0
M7 2 3 10 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=24470 $Y=110705 $dt=0
M8 17 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=25710 $Y=76905 $dt=0
M9 15 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=25710 $Y=110705 $dt=0
M10 2 3 16 2 ne3i L=4e-07 W=3e-05 AD=3.39e-11 AS=1.5e-13 PD=3.226e-05 PS=6.001e-05 $X=33470 $Y=76905 $dt=0
M11 2 3 14 2 ne3i L=4e-07 W=3e-05 AD=3.39e-11 AS=1.5e-13 PD=3.226e-05 PS=6.001e-05 $X=33470 $Y=110705 $dt=0
M12 20 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=3.39e-11 PD=6.001e-05 PS=3.226e-05 $X=36130 $Y=76905 $dt=0
M13 18 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=3.39e-11 PD=6.001e-05 PS=3.226e-05 $X=36130 $Y=110705 $dt=0
M14 2 3 21 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=43890 $Y=76905 $dt=0
M15 2 3 19 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=43890 $Y=110705 $dt=0
M16 24 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=45130 $Y=76905 $dt=0
M17 22 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=45130 $Y=110705 $dt=0
M18 2 3 25 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=52890 $Y=76905 $dt=0
M19 2 3 23 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=52890 $Y=110705 $dt=0
M20 28 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=54130 $Y=76905 $dt=0
M21 26 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=54130 $Y=110705 $dt=0
M22 2 3 29 2 ne3i L=4e-07 W=3e-05 AD=1.89e-11 AS=1.5e-13 PD=6.126e-05 PS=6.001e-05 $X=61890 $Y=76905 $dt=0
M23 2 3 27 2 ne3i L=4e-07 W=3e-05 AD=1.89e-11 AS=1.5e-13 PD=6.126e-05 PS=6.001e-05 $X=61890 $Y=110705 $dt=0
D24 5 1 ddnwmv AREA=4.69976e-09 PJ=0.00027464 perimeter=0.00027464 $X=2570 $Y=72575 $dt=2
D25 2 1 dipdnwmv AREA=4.16648e-09 PJ=0.00025864 perimeter=0.00025864 $X=4570 $Y=74575 $dt=4
.ends jio_base_ntrc_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_basepsc_pc                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_basepsc_pc 1 2 3 4
** N=42 EP=4 FDC=149
X1073 2 3 18 17 jio_pe3isb_pc $T=14365 150990 1 180 $X=6700 $Y=149060
X1074 2 3 16 15 jio_pe3isb_pc $T=14365 184790 1 180 $X=6700 $Y=182860
X1075 2 3 14 13 jio_pe3isb_pc $T=20965 150990 1 180 $X=13300 $Y=149060
X1076 2 3 12 11 jio_pe3isb_pc $T=20965 184790 1 180 $X=13300 $Y=182860
X1077 2 3 26 25 jio_pe3isb_pc $T=27565 150990 1 180 $X=19900 $Y=149060
X1078 2 3 24 23 jio_pe3isb_pc $T=27565 184790 1 180 $X=19900 $Y=182860
X1079 2 3 22 21 jio_pe3isb_pc $T=34165 150990 1 180 $X=26500 $Y=149060
X1080 2 3 20 19 jio_pe3isb_pc $T=34165 184790 1 180 $X=26500 $Y=182860
X1081 2 3 34 33 jio_pe3isb_pc $T=35835 150990 0 0 $X=35120 $Y=149060
X1082 2 3 32 31 jio_pe3isb_pc $T=35835 184790 0 0 $X=35120 $Y=182860
X1083 2 3 30 29 jio_pe3isb_pc $T=42435 150990 0 0 $X=41720 $Y=149060
X1084 2 3 28 27 jio_pe3isb_pc $T=42435 184790 0 0 $X=41720 $Y=182860
X1085 2 3 42 41 jio_pe3isb_pc $T=49035 150990 0 0 $X=48320 $Y=149060
X1086 2 3 40 39 jio_pe3isb_pc $T=49035 184790 0 0 $X=48320 $Y=182860
X1087 2 3 38 37 jio_pe3isb_pc $T=55635 150990 0 0 $X=54920 $Y=149060
X1088 2 3 36 35 jio_pe3isb_pc $T=55635 184790 0 0 $X=54920 $Y=182860
X1276 2 4 10 3 1 jio_base_ntrc_pc $T=0 0 0 0 $X=2560 $Y=72565
M0 18 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=8060 $Y=152815 $dt=1
M1 16 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=8060 $Y=186615 $dt=1
M2 2 9 17 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=13370 $Y=152815 $dt=1
M3 2 9 15 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=13370 $Y=186615 $dt=1
M4 14 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=14660 $Y=152815 $dt=1
M5 12 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=14660 $Y=186615 $dt=1
M6 2 9 13 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=19970 $Y=152815 $dt=1
M7 2 9 11 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=19970 $Y=186615 $dt=1
M8 26 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=21260 $Y=152815 $dt=1
M9 24 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=21260 $Y=186615 $dt=1
M10 2 9 25 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=26570 $Y=152815 $dt=1
M11 2 9 23 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=26570 $Y=186615 $dt=1
M12 22 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=27860 $Y=152815 $dt=1
M13 20 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=27860 $Y=186615 $dt=1
M14 2 9 21 2 pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=33170 $Y=152815 $dt=1
M15 2 9 19 2 pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=33170 $Y=186615 $dt=1
M16 33 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=36480 $Y=152815 $dt=1
M17 31 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=36480 $Y=186615 $dt=1
M18 2 9 34 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=41790 $Y=152815 $dt=1
M19 2 9 32 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=41790 $Y=186615 $dt=1
M20 29 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=43080 $Y=152815 $dt=1
M21 27 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=43080 $Y=186615 $dt=1
M22 2 9 30 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=48390 $Y=152815 $dt=1
M23 2 9 28 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=48390 $Y=186615 $dt=1
M24 41 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=49680 $Y=152815 $dt=1
M25 39 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=49680 $Y=186615 $dt=1
M26 2 9 42 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=54990 $Y=152815 $dt=1
M27 2 9 40 2 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=54990 $Y=186615 $dt=1
M28 37 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=56280 $Y=152815 $dt=1
M29 35 9 2 2 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=56280 $Y=186615 $dt=1
M30 2 9 38 2 pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=61590 $Y=152815 $dt=1
M31 2 9 36 2 pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=61590 $Y=186615 $dt=1
D32 1 2 p_ddnwmv AREA=4.5084e-09 PJ=0.00026872 perimeter=0.00026872 $X=2500 $Y=150035 $dt=3
R33 9 2 L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=2 $X=4475 $Y=153720 $dt=7
R34 10 4 L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=2 $X=65085 $Y=153720 $dt=7
D35 9 2 p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=4475 $Y=152700 $dt=12
D36 2 2 p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=4475 $Y=157020 $dt=12
D37 10 2 p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=65085 $Y=152700 $dt=12
D38 4 2 p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=65085 $Y=157020 $dt=12
.ends jio_basepsc_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VDDPADPC                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VDDPADPC VDD3I GNDI VDDRI VDDOI GNDRI GNDOI PSUB
** N=7 EP=7 FDC=149
X0 PSUB VDDOI VDD3I GNDOI jio_basepsc_pc $T=0 0 0 0 $X=-320 $Y=0
.ends VDDPADPC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_base_ptrpsfl_pc                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_base_ptrpsfl_pc 1 3
** N=3 EP=2 FDC=17
D0 3 1 p_ddnwmv AREA=4.5084e-09 PJ=0.00026872 perimeter=0.00026872 $X=2500 $Y=150035 $dt=3
D1 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=13480 $Y=153600 $dt=12
D2 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=13480 $Y=187400 $dt=12
D3 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=20080 $Y=153600 $dt=12
D4 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=20080 $Y=187400 $dt=12
D5 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=26680 $Y=153600 $dt=12
D6 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=26680 $Y=187400 $dt=12
D7 1 1 p_dp3 AREA=3.4348e-11 PJ=3.018e-05 perimeter=3.018e-05 $X=33280 $Y=153600 $dt=12
D8 1 1 p_dp3 AREA=3.4348e-11 PJ=3.018e-05 perimeter=3.018e-05 $X=33280 $Y=187400 $dt=12
D9 1 1 p_dp3 AREA=3.4348e-11 PJ=3.018e-05 perimeter=3.018e-05 $X=35480 $Y=153600 $dt=12
D10 1 1 p_dp3 AREA=3.4348e-11 PJ=3.018e-05 perimeter=3.018e-05 $X=35480 $Y=187400 $dt=12
D11 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=41900 $Y=153600 $dt=12
D12 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=41900 $Y=187400 $dt=12
D13 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=48500 $Y=153600 $dt=12
D14 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=48500 $Y=187400 $dt=12
D15 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=55100 $Y=153600 $dt=12
D16 1 1 p_dp3 AREA=3.9334e-11 PJ=5.824e-05 perimeter=5.824e-05 $X=55100 $Y=187400 $dt=12
.ends jio_base_ptrpsfl_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_base_ntr_pc                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_base_ntr_pc 1 2 3 4 5 6 7
** N=31 EP=7 FDC=62
X100 2 6 10 11 jio_ne3isb_pc $T=16420 75080 1 180 $X=6100 $Y=73130
X101 2 6 8 9 jio_ne3isb_pc $T=16420 108880 1 180 $X=6100 $Y=106930
X102 2 6 14 15 jio_ne3isb_pc $T=25420 75080 1 180 $X=15100 $Y=73130
X103 2 6 12 13 jio_ne3isb_pc $T=25420 108880 1 180 $X=15100 $Y=106930
X104 2 6 18 19 jio_ne3isb_pc $T=34420 75080 1 180 $X=24100 $Y=73130
X105 2 6 16 17 jio_ne3isb_pc $T=34420 108880 1 180 $X=24100 $Y=106930
X106 2 6 22 23 jio_ne3isb_pc $T=35580 75080 0 0 $X=34520 $Y=73130
X107 2 6 20 21 jio_ne3isb_pc $T=35580 108880 0 0 $X=34520 $Y=106930
X108 2 6 26 27 jio_ne3isb_pc $T=44580 75080 0 0 $X=43520 $Y=73130
X109 2 6 24 25 jio_ne3isb_pc $T=44580 108880 0 0 $X=43520 $Y=106930
X110 2 6 30 31 jio_ne3isb_pc $T=53580 75080 0 0 $X=52520 $Y=73130
X111 2 6 28 29 jio_ne3isb_pc $T=53580 108880 0 0 $X=52520 $Y=106930
M0 11 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.89e-11 PD=6.001e-05 PS=6.126e-05 $X=7710 $Y=76905 $dt=0
M1 9 4 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.89e-11 PD=6.001e-05 PS=6.126e-05 $X=7710 $Y=110705 $dt=0
M2 2 3 10 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=15470 $Y=76905 $dt=0
M3 2 3 8 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=15470 $Y=110705 $dt=0
M4 15 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=16710 $Y=76905 $dt=0
M5 13 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=16710 $Y=110705 $dt=0
M6 2 3 14 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=24470 $Y=76905 $dt=0
M7 2 3 12 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=24470 $Y=110705 $dt=0
M8 19 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=25710 $Y=76905 $dt=0
M9 17 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=25710 $Y=110705 $dt=0
M10 2 3 18 2 ne3i L=4e-07 W=3e-05 AD=3.39e-11 AS=1.5e-13 PD=3.226e-05 PS=6.001e-05 $X=33470 $Y=76905 $dt=0
M11 2 3 16 2 ne3i L=4e-07 W=3e-05 AD=3.39e-11 AS=1.5e-13 PD=3.226e-05 PS=6.001e-05 $X=33470 $Y=110705 $dt=0
M12 22 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=3.39e-11 PD=6.001e-05 PS=3.226e-05 $X=36130 $Y=76905 $dt=0
M13 20 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=3.39e-11 PD=6.001e-05 PS=3.226e-05 $X=36130 $Y=110705 $dt=0
M14 2 3 23 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=43890 $Y=76905 $dt=0
M15 2 3 21 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=43890 $Y=110705 $dt=0
M16 26 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=45130 $Y=76905 $dt=0
M17 24 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=45130 $Y=110705 $dt=0
M18 2 3 27 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=52890 $Y=76905 $dt=0
M19 2 3 25 2 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=52890 $Y=110705 $dt=0
M20 30 3 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=54130 $Y=76905 $dt=0
M21 28 5 2 2 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=54130 $Y=110705 $dt=0
M22 2 3 31 2 ne3i L=4e-07 W=3e-05 AD=1.89e-11 AS=1.5e-13 PD=6.126e-05 PS=6.001e-05 $X=61890 $Y=76905 $dt=0
M23 2 5 29 2 ne3i L=4e-07 W=3e-05 AD=1.89e-11 AS=1.5e-13 PD=6.126e-05 PS=6.001e-05 $X=61890 $Y=110705 $dt=0
D24 7 1 ddnwmv AREA=4.69976e-09 PJ=0.00027464 perimeter=0.00027464 $X=2570 $Y=72575 $dt=2
D25 2 1 dipdnwmv AREA=4.16648e-09 PJ=0.00025864 perimeter=0.00025864 $X=4570 $Y=74575 $dt=4
.ends jio_base_ntr_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VDDORPADPC                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VDDORPADPC PSUB VDDORI GNDOI VDD3I GNDI GNDRI
** N=7 EP=6 FDC=82
X1219 VDDORI PSUB jio_base_ptrpsfl_pc $T=0 0 0 0 $X=510 $Y=137985
X1220 VDDORI GNDOI 7 7 7 VDDORI PSUB jio_base_ntr_pc $T=0 0 0 0 $X=2560 $Y=72565
R0 7 GNDOI L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=VDDORI $X=65085 $Y=153720 $dt=7
D1 7 VDDORI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=65085 $Y=152700 $dt=12
D2 GNDOI VDDORI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=65085 $Y=157020 $dt=12
.ends VDDORPADPC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: GNDPADPC                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt GNDPADPC GNDI VDD3I VDDRI VDDOI GNDRI GNDOI PSUB
** N=7 EP=7 FDC=149
X0 PSUB VDDOI GNDI GNDOI jio_basepsc_pc $T=0 0 0 0 $X=-320 $Y=0
.ends GNDPADPC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: GNDORPADPC                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt GNDORPADPC PSUB VDDOI GNDORI VDD3I GNDI VDDRI
** N=31 EP=6 FDC=66
X1949 GNDORI VDDOI 10 11 jio_ne3isbg_pc $T=16420 150990 1 180 $X=6100 $Y=149915
X1950 GNDORI VDDOI 8 9 jio_ne3isbg_pc $T=16420 184790 1 180 $X=6100 $Y=183715
X1951 GNDORI VDDOI 14 15 jio_ne3isbg_pc $T=25420 150990 1 180 $X=15100 $Y=149915
X1952 GNDORI VDDOI 12 13 jio_ne3isbg_pc $T=25420 184790 1 180 $X=15100 $Y=183715
X1953 GNDORI VDDOI 22 23 jio_ne3isbg_pc $T=34420 150990 1 180 $X=24100 $Y=149915
X1954 GNDORI VDDOI 20 21 jio_ne3isbg_pc $T=34420 184790 1 180 $X=24100 $Y=183715
X1955 GNDORI VDDOI 18 19 jio_ne3isbg_pc $T=35580 150990 0 0 $X=34520 $Y=149915
X1956 GNDORI VDDOI 16 17 jio_ne3isbg_pc $T=35580 184790 0 0 $X=34520 $Y=183715
X1957 GNDORI VDDOI 26 27 jio_ne3isbg_pc $T=44580 150990 0 0 $X=43520 $Y=149915
X1958 GNDORI VDDOI 24 25 jio_ne3isbg_pc $T=44580 184790 0 0 $X=43520 $Y=183715
X1959 GNDORI VDDOI 30 31 jio_ne3isbg_pc $T=53580 150990 0 0 $X=52520 $Y=149915
X1960 GNDORI VDDOI 28 29 jio_ne3isbg_pc $T=53580 184790 0 0 $X=52520 $Y=183715
M0 11 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.89e-11 PD=6.001e-05 PS=6.126e-05 $X=7710 $Y=152815 $dt=0
M1 9 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.89e-11 PD=6.001e-05 PS=6.126e-05 $X=7710 $Y=186615 $dt=0
M2 GNDORI 7 10 GNDORI ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=15470 $Y=152815 $dt=0
M3 GNDORI 7 8 GNDORI ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=15470 $Y=186615 $dt=0
M4 15 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=16710 $Y=152815 $dt=0
M5 13 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=16710 $Y=186615 $dt=0
M6 GNDORI 7 14 GNDORI ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=24470 $Y=152815 $dt=0
M7 GNDORI 7 12 GNDORI ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=24470 $Y=186615 $dt=0
M8 23 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=25710 $Y=152815 $dt=0
M9 21 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=25710 $Y=186615 $dt=0
M10 GNDORI 7 22 GNDORI ne3i L=4e-07 W=3e-05 AD=3.39e-11 AS=1.5e-13 PD=3.226e-05 PS=6.001e-05 $X=33470 $Y=152815 $dt=0
M11 GNDORI 7 20 GNDORI ne3i L=4e-07 W=3e-05 AD=3.39e-11 AS=1.5e-13 PD=3.226e-05 PS=6.001e-05 $X=33470 $Y=186615 $dt=0
M12 18 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=3.39e-11 PD=6.001e-05 PS=3.226e-05 $X=36130 $Y=152815 $dt=0
M13 16 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=3.39e-11 PD=6.001e-05 PS=3.226e-05 $X=36130 $Y=186615 $dt=0
M14 GNDORI 7 19 GNDORI ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=43890 $Y=152815 $dt=0
M15 GNDORI 7 17 GNDORI ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=43890 $Y=186615 $dt=0
M16 26 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=45130 $Y=152815 $dt=0
M17 24 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=45130 $Y=186615 $dt=0
M18 GNDORI 7 27 GNDORI ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=52890 $Y=152815 $dt=0
M19 GNDORI 7 25 GNDORI ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=52890 $Y=186615 $dt=0
M20 30 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=54130 $Y=152815 $dt=0
M21 28 7 GNDORI GNDORI ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=54130 $Y=186615 $dt=0
M22 GNDORI 7 31 GNDORI ne3i L=4e-07 W=3e-05 AD=1.89e-11 AS=1.5e-13 PD=6.126e-05 PS=6.001e-05 $X=61890 $Y=152815 $dt=0
M23 GNDORI 7 29 GNDORI ne3i L=4e-07 W=3e-05 AD=1.89e-11 AS=1.5e-13 PD=6.126e-05 PS=6.001e-05 $X=61890 $Y=186615 $dt=0
D24 PSUB VDDOI ddnwmv AREA=4.69976e-09 PJ=0.00027464 perimeter=0.00027464 $X=2570 $Y=148485 $dt=2
D25 GNDORI VDDOI dipdnwmv AREA=4.16648e-09 PJ=0.00025864 perimeter=0.00025864 $X=4570 $Y=150485 $dt=4
R26 GNDORI 7 L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=VDDOI $X=4810 $Y=136135 $dt=6
D27 GNDORI VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=4810 $Y=135115 $dt=11
D28 7 VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=4810 $Y=139435 $dt=11
D29 PSUB VDDOI p_dnw3 AREA=4.54356e-09 PJ=0.00026992 perimeter=0.00026992 $X=2840 $Y=72575 $dt=13
.ends GNDORPADPC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_base_ptr_pc                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_base_ptr_pc 1 2 3 4 5 6 7
** N=31 EP=7 FDC=63
X37 1 3 9 8 jio_pe3isb_pc $T=14365 150990 1 180 $X=6700 $Y=149060
X38 1 3 11 10 jio_pe3isb_pc $T=20965 150990 1 180 $X=13300 $Y=149060
X39 1 3 19 18 jio_pe3isb_pc $T=27565 150990 1 180 $X=19900 $Y=149060
X40 1 3 17 16 jio_pe3isb_pc $T=27565 184790 1 180 $X=19900 $Y=182860
X41 1 3 15 14 jio_pe3isb_pc $T=34165 150990 1 180 $X=26500 $Y=149060
X42 1 3 13 12 jio_pe3isb_pc $T=34165 184790 1 180 $X=26500 $Y=182860
X43 1 3 27 26 jio_pe3isb_pc $T=35835 150990 0 0 $X=35120 $Y=149060
X44 1 3 25 24 jio_pe3isb_pc $T=35835 184790 0 0 $X=35120 $Y=182860
X45 1 3 23 22 jio_pe3isb_pc $T=42435 150990 0 0 $X=41720 $Y=149060
X46 1 3 21 20 jio_pe3isb_pc $T=42435 184790 0 0 $X=41720 $Y=182860
X47 1 3 29 28 jio_pe3isb_pc $T=49035 150990 0 0 $X=48320 $Y=149060
X48 1 3 31 30 jio_pe3isb_pc $T=55635 150990 0 0 $X=54920 $Y=149060
M0 9 4 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=8060 $Y=152815 $dt=1
M1 1 4 8 1 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=13370 $Y=152815 $dt=1
M2 11 4 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=14660 $Y=152815 $dt=1
M3 1 4 10 1 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=19970 $Y=152815 $dt=1
M4 19 4 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=21260 $Y=152815 $dt=1
M5 17 5 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=21260 $Y=186615 $dt=1
M6 1 4 18 1 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=26570 $Y=152815 $dt=1
M7 1 5 16 1 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=26570 $Y=186615 $dt=1
M8 15 4 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=27860 $Y=152815 $dt=1
M9 13 5 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=27860 $Y=186615 $dt=1
M10 1 4 14 1 pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=33170 $Y=152815 $dt=1
M11 1 4 12 1 pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=33170 $Y=186615 $dt=1
M12 26 4 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=36480 $Y=152815 $dt=1
M13 24 4 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=36480 $Y=186615 $dt=1
M14 1 4 27 1 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=41790 $Y=152815 $dt=1
M15 1 4 25 1 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=41790 $Y=186615 $dt=1
M16 22 4 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=43080 $Y=152815 $dt=1
M17 20 4 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=43080 $Y=186615 $dt=1
M18 1 4 23 1 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=48390 $Y=152815 $dt=1
M19 1 4 21 1 pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=48390 $Y=186615 $dt=1
M20 28 4 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=49680 $Y=152815 $dt=1
M21 1 6 29 1 pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=54990 $Y=152815 $dt=1
M22 30 6 1 1 pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=56280 $Y=152815 $dt=1
M23 1 6 31 1 pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=61590 $Y=152815 $dt=1
D24 7 1 p_ddnwmv AREA=4.5084e-09 PJ=0.00026872 perimeter=0.00026872 $X=2500 $Y=150035 $dt=3
D25 2 1 dipdnwmv AREA=2.1664e-10 PJ=5.908e-05 perimeter=5.908e-05 $X=4500 $Y=201395 $dt=4
D26 2 1 dipdnwmv AREA=2.1664e-10 PJ=5.908e-05 perimeter=5.908e-05 $X=51960 $Y=201395 $dt=4
.ends jio_base_ptr_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_baseti_pc                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_baseti_pc 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14
** N=14 EP=14 FDC=131
X61 2 5 13 14 12 8 1 jio_base_ntr_pc $T=0 0 0 0 $X=2560 $Y=72565
X62 2 5 8 9 11 10 1 jio_base_ptr_pc $T=0 0 0 0 $X=2500 $Y=149060
D0 1 2 ddnwmv AREA=5.2955e-10 PJ=0.00010026 perimeter=0.00010026 $X=2500 $Y=224395 $dt=2
D1 1 6 ddnwmv AREA=3.7825e-10 PJ=8.026e-05 perimeter=8.026e-05 $X=42500 $Y=224395 $dt=2
D2 1 3 p_ddnwmv AREA=9.789e-10 PJ=0.00016012 perimeter=0.00016012 $X=2500 $Y=244525 $dt=3
D3 5 2 dipdnwmv AREA=1.9592e-10 PJ=7.464e-05 perimeter=7.464e-05 $X=4500 $Y=226395 $dt=4
D4 4 3 dipdnwmv AREA=3.1903e-10 PJ=0.00013246 perimeter=0.00013246 $X=4500 $Y=246525 $dt=4
D5 7 6 dipdnwmv AREA=1.3272e-10 PJ=5.464e-05 perimeter=5.464e-05 $X=44500 $Y=226395 $dt=4
.ends jio_baseti_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ICPC                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ICPC VDDOI VDD3I PSUB GNDI GNDOI VDDRI GNDRI Y PAD PO
+ PI
** N=26 EP=11 FDC=190
X415 PSUB VDDOI VDD3I GNDI GNDOI VDDRI GNDRI PAD 12 12
+ 12 15 15 15 jio_baseti_pc $T=0 0 0 0 $X=-320 $Y=0
M0 15 12 GNDOI GNDOI ne3i L=4e-07 W=1.2e-06 AD=6.36e-13 AS=6.36e-13 PD=3.46e-06 PS=3.46e-06 $X=10900 $Y=214545 $dt=0
M1 GNDI 22 14 GNDI ne3i L=4e-07 W=1.2e-06 AD=4.02e-13 AS=6.12e-13 PD=1.87e-06 PS=3.42e-06 $X=43225 $Y=248510 $dt=0
M2 14 22 GNDI GNDI ne3i L=4e-07 W=1.2e-06 AD=6.24e-13 AS=4.02e-13 PD=3.44e-06 PS=1.87e-06 $X=44295 $Y=248510 $dt=0
M3 16 14 GNDI GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=8.064e-13 PD=2.22e-06 PS=4.32e-06 $X=48745 $Y=248340 $dt=0
M4 GNDI 14 16 GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=4.536e-13 PD=2.22e-06 PS=2.22e-06 $X=49685 $Y=248340 $dt=0
M5 16 14 GNDI GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=4.536e-13 PD=2.22e-06 PS=2.22e-06 $X=50625 $Y=248340 $dt=0
M6 GNDI 14 16 GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=4.536e-13 PD=2.22e-06 PS=2.22e-06 $X=51565 $Y=248340 $dt=0
M7 17 14 GNDI GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=4.536e-13 PD=2.22e-06 PS=2.22e-06 $X=52505 $Y=248340 $dt=0
M8 GNDI 14 17 GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=4.536e-13 PD=2.22e-06 PS=2.22e-06 $X=53445 $Y=248340 $dt=0
M9 19 GNDOI GNDOI GNDOI ne3i L=4e-07 W=1.2e-05 AD=6e-14 AS=6.66e-12 PD=2.401e-05 PS=2.511e-05 $X=53865 $Y=203375 $dt=0
M10 Y 16 GNDI GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=4.536e-13 PD=2.22e-06 PS=2.22e-06 $X=54385 $Y=248340 $dt=0
M11 GNDI 16 Y GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=4.536e-13 PD=2.22e-06 PS=2.22e-06 $X=55325 $Y=248340 $dt=0
M12 GNDRI 20 22 GNDRI ne3i L=4e-07 W=2e-06 AD=5.4e-13 AS=9.6e-13 PD=2.54e-06 PS=4.96e-06 $X=55490 $Y=228495 $dt=0
M13 Y 16 GNDI GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=4.536e-13 PD=2.22e-06 PS=2.22e-06 $X=56265 $Y=248340 $dt=0
M14 22 20 GNDRI GNDRI ne3i L=4e-07 W=2e-06 AD=5.4e-13 AS=5.4e-13 PD=2.54e-06 PS=2.54e-06 $X=56430 $Y=228495 $dt=0
M15 GNDI 16 Y GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=4.536e-13 PD=2.22e-06 PS=2.22e-06 $X=57205 $Y=248340 $dt=0
M16 GNDRI 20 22 GNDRI ne3i L=4e-07 W=2e-06 AD=9.6e-13 AS=5.4e-13 PD=4.96e-06 PS=2.54e-06 $X=57370 $Y=228495 $dt=0
M17 GNDOI GNDOI 21 GNDOI ne3i L=4e-07 W=1.2e-05 AD=6.66e-12 AS=6e-14 PD=2.511e-05 PS=2.401e-05 $X=57565 $Y=203375 $dt=0
M18 Y 16 GNDI GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=4.536e-13 PD=2.22e-06 PS=2.22e-06 $X=58145 $Y=248340 $dt=0
M19 GNDI 16 Y GNDI ne3i L=4e-07 W=1.68e-06 AD=8.064e-13 AS=4.536e-13 PD=4.32e-06 PS=2.22e-06 $X=59085 $Y=248340 $dt=0
M20 18 14 PO GNDI ne3i L=4e-07 W=1.68e-06 AD=4.536e-13 AS=8.064e-13 PD=2.22e-06 PS=4.32e-06 $X=62265 $Y=248110 $dt=0
M21 GNDI PI 18 GNDI ne3i L=4e-07 W=1.68e-06 AD=8.064e-13 AS=4.536e-13 PD=4.32e-06 PS=2.22e-06 $X=63205 $Y=248110 $dt=0
M22 20 VDDOI VDDOI VDDOI pe3i L=3.5e-07 W=1.2e-05 AD=6.78e-12 AS=6.24e-12 PD=1.313e-05 PS=2.504e-05 $X=22325 $Y=234735 $dt=1
M23 VDDOI VDDOI 20 VDDOI pe3i L=3.5e-07 W=1.2e-05 AD=6.24e-12 AS=6.78e-12 PD=2.504e-05 PS=1.313e-05 $X=22325 $Y=236215 $dt=1
M24 14 22 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=1.152e-12 PD=2.94e-06 PS=5.76e-06 $X=42235 $Y=254765 $dt=1
M25 VDD3I 22 14 VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=1.152e-12 AS=6.48e-13 PD=5.76e-06 PS=2.94e-06 $X=43125 $Y=254765 $dt=1
M26 16 14 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=1.152e-12 PD=2.94e-06 PS=5.76e-06 $X=45125 $Y=254765 $dt=1
M27 VDD3I 14 16 VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=46015 $Y=254765 $dt=1
M28 17 14 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=46905 $Y=254765 $dt=1
M29 VDD3I 14 17 VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=47795 $Y=254765 $dt=1
M30 17 14 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=48685 $Y=254765 $dt=1
M31 VDD3I 14 17 VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=49575 $Y=254765 $dt=1
M32 17 14 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=50465 $Y=254765 $dt=1
M33 VDD3I 14 17 VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=51355 $Y=254765 $dt=1
M34 Y 17 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=52245 $Y=254765 $dt=1
M35 VDD3I 17 Y VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=53135 $Y=254765 $dt=1
M36 Y 17 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=54025 $Y=254765 $dt=1
M37 VDD3I 17 Y VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=54915 $Y=254765 $dt=1
M38 22 20 VDDRI VDDRI pe3i L=3.5e-07 W=2.2e-06 AD=6.49e-13 AS=1.111e-12 PD=2.79e-06 PS=5.41e-06 $X=55515 $Y=234765 $dt=1
M39 Y 17 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=55805 $Y=254765 $dt=1
M40 VDDRI 20 22 VDDRI pe3i L=3.5e-07 W=2.2e-06 AD=6.49e-13 AS=6.49e-13 PD=2.79e-06 PS=2.79e-06 $X=56455 $Y=234765 $dt=1
M41 VDD3I 17 Y VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=56695 $Y=254765 $dt=1
M42 22 20 VDDRI VDDRI pe3i L=3.5e-07 W=2.2e-06 AD=6.49e-13 AS=6.49e-13 PD=2.79e-06 PS=2.79e-06 $X=57395 $Y=234765 $dt=1
M43 Y 17 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=57585 $Y=254765 $dt=1
M44 VDDRI 20 22 VDDRI pe3i L=3.5e-07 W=2.2e-06 AD=6.49e-13 AS=6.49e-13 PD=2.79e-06 PS=2.79e-06 $X=58335 $Y=234765 $dt=1
M45 VDD3I 17 Y VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=58475 $Y=254765 $dt=1
M46 22 20 VDDRI VDDRI pe3i L=3.5e-07 W=2.2e-06 AD=6.49e-13 AS=6.49e-13 PD=2.79e-06 PS=2.79e-06 $X=59275 $Y=234765 $dt=1
M47 Y 17 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=6.48e-13 PD=2.94e-06 PS=2.94e-06 $X=59365 $Y=254765 $dt=1
M48 VDDRI 20 22 VDDRI pe3i L=3.5e-07 W=2.2e-06 AD=1.111e-12 AS=6.49e-13 PD=5.41e-06 PS=2.79e-06 $X=60215 $Y=234765 $dt=1
M49 VDD3I 17 Y VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=1.152e-12 AS=6.48e-13 PD=5.76e-06 PS=2.94e-06 $X=60255 $Y=254765 $dt=1
M50 PO 14 VDD3I VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=6.48e-13 AS=1.248e-12 PD=2.94e-06 PS=5.84e-06 $X=62365 $Y=254765 $dt=1
M51 VDD3I PI PO VDD3I pe3i L=3.5e-07 W=2.4e-06 AD=1.152e-12 AS=6.48e-13 PD=5.76e-06 PS=2.94e-06 $X=63255 $Y=254765 $dt=1
R52 19 20 L=1.32e-06 W=1.2e-05 $[rdn3] $SUB=GNDOI $X=54270 $Y=203375 $dt=5
R53 20 21 L=1.32e-06 W=1.2e-05 $[rdn3] $SUB=GNDOI $X=56245 $Y=203375 $dt=5
R54 VDDOI 12 L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=VDDOI $X=3990 $Y=178955 $dt=7
D55 GNDOI 20 dn3 AREA=7.92e-12 PJ=1.32e-06 perimeter=1.32e-06 $X=55585 $Y=203375 $dt=9
D56 VDDOI VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=3990 $Y=177935 $dt=12
D57 12 VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=3990 $Y=182255 $dt=12
R58 20 PAD L=4.5e-06 W=2.5e-06 $[rpp1] $X=52790 $Y=196775 $dt=14
.ends ICPC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BT4PC                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BT4PC VDD3I VDDOI GNDOI A PSUB GNDI EN VDDRI GNDRI PAD
** N=27 EP=10 FDC=183
X421 PSUB VDDOI VDD3I GNDI GNDOI VDDRI GNDRI PAD 11 21
+ 22 23 19 15 jio_baseti_pc $T=0 0 0 0 $X=-320 $Y=0
M0 15 16 GNDOI GNDOI ne3i L=4e-07 W=5.5e-06 AD=1.76e-12 AS=2.915e-12 PD=6.14e-06 PS=1.206e-05 $X=6380 $Y=203055 $dt=0
M1 18 EN GNDI GNDI ne3i L=4e-07 W=1.1e-06 AD=5.28e-13 AS=5.28e-13 PD=3.16e-06 PS=3.16e-06 $X=6395 $Y=248525 $dt=0
M2 GNDOI 16 15 GNDOI ne3i L=4e-07 W=5.5e-06 AD=2.915e-12 AS=1.76e-12 PD=1.206e-05 PS=6.14e-06 $X=7420 $Y=203055 $dt=0
M3 GNDI A 24 GNDI ne3i L=4e-07 W=1.1e-06 AD=2.97e-13 AS=5.28e-13 PD=1.64e-06 PS=3.16e-06 $X=8035 $Y=248525 $dt=0
M4 14 17 GNDOI GNDOI ne3i L=4e-07 W=1.3e-06 AD=3.51e-13 AS=6.24e-13 PD=1.84e-06 PS=3.56e-06 $X=8915 $Y=228445 $dt=0
M5 24 A GNDI GNDI ne3i L=4e-07 W=1.1e-06 AD=2.97e-13 AS=2.97e-13 PD=1.64e-06 PS=1.64e-06 $X=8975 $Y=248525 $dt=0
M6 22 14 GNDOI GNDOI ne3i L=4e-07 W=6.1e-06 AD=3.233e-12 AS=3.233e-12 PD=1.326e-05 PS=1.326e-05 $X=9160 $Y=209645 $dt=0
M7 GNDOI 17 14 GNDOI ne3i L=4e-07 W=1.3e-06 AD=3.51e-13 AS=3.51e-13 PD=1.84e-06 PS=1.84e-06 $X=9855 $Y=228445 $dt=0
M8 17 18 24 GNDI ne3i L=4e-07 W=1.1e-06 AD=2.97e-13 AS=2.97e-13 PD=1.64e-06 PS=1.64e-06 $X=9915 $Y=248525 $dt=0
M9 14 17 GNDOI GNDOI ne3i L=4e-07 W=1.3e-06 AD=3.51e-13 AS=3.51e-13 PD=1.84e-06 PS=1.84e-06 $X=10795 $Y=228445 $dt=0
M10 24 18 17 GNDI ne3i L=4e-07 W=1.1e-06 AD=5.28e-13 AS=2.97e-13 PD=3.16e-06 PS=1.64e-06 $X=10855 $Y=248525 $dt=0
M11 19 11 GNDOI GNDOI ne3i L=4e-07 W=1.2e-06 AD=6.36e-13 AS=6.36e-13 PD=3.46e-06 PS=3.46e-06 $X=10900 $Y=212165 $dt=0
M12 GNDOI 17 14 GNDOI ne3i L=4e-07 W=1.3e-06 AD=3.51e-13 AS=3.51e-13 PD=1.84e-06 PS=1.84e-06 $X=11735 $Y=228445 $dt=0
M13 16 20 GNDOI GNDOI ne3i L=4e-07 W=1.3e-06 AD=3.51e-13 AS=3.51e-13 PD=1.84e-06 PS=1.84e-06 $X=12675 $Y=228445 $dt=0
M14 20 A GNDI GNDI ne3i L=4e-07 W=1.1e-06 AD=2.97e-13 AS=5.28e-13 PD=1.64e-06 PS=3.16e-06 $X=13535 $Y=248525 $dt=0
M15 GNDOI 20 16 GNDOI ne3i L=4e-07 W=1.3e-06 AD=3.51e-13 AS=3.51e-13 PD=1.84e-06 PS=1.84e-06 $X=13615 $Y=228445 $dt=0
M16 GNDI A 20 GNDI ne3i L=4e-07 W=1.1e-06 AD=2.97e-13 AS=2.97e-13 PD=1.64e-06 PS=1.64e-06 $X=14475 $Y=248525 $dt=0
M17 16 20 GNDOI GNDOI ne3i L=4e-07 W=1.3e-06 AD=3.51e-13 AS=3.51e-13 PD=1.84e-06 PS=1.84e-06 $X=14555 $Y=228445 $dt=0
M18 20 EN GNDI GNDI ne3i L=4e-07 W=1.1e-06 AD=2.97e-13 AS=2.97e-13 PD=1.64e-06 PS=1.64e-06 $X=15415 $Y=248525 $dt=0
M19 GNDOI 20 16 GNDOI ne3i L=4e-07 W=1.3e-06 AD=6.24e-13 AS=3.51e-13 PD=3.56e-06 PS=1.84e-06 $X=15495 $Y=228445 $dt=0
M20 GNDI EN 20 GNDI ne3i L=4e-07 W=1.1e-06 AD=5.28e-13 AS=2.97e-13 PD=3.16e-06 PS=1.64e-06 $X=16355 $Y=248525 $dt=0
M21 25 14 21 GNDOI ne3i L=4e-07 W=3.7e-06 AD=1.961e-12 AS=1.961e-12 PD=8.46e-06 PS=8.46e-06 $X=60440 $Y=207685 $dt=0
M22 25 14 GNDOI GNDOI ne3i L=4e-07 W=3.7e-06 AD=1.961e-12 AS=1.961e-12 PD=8.46e-06 PS=8.46e-06 $X=60440 $Y=212045 $dt=0
M23 23 16 GNDOI GNDOI ne3i L=4e-07 W=8e-06 AD=2.56e-12 AS=4.24e-12 PD=8.64e-06 PS=1.706e-05 $X=62180 $Y=207745 $dt=0
M24 GNDOI 16 23 GNDOI ne3i L=4e-07 W=8e-06 AD=4.24e-12 AS=2.56e-12 PD=1.706e-05 PS=8.64e-06 $X=63220 $Y=207745 $dt=0
M25 15 16 VDDOI VDDOI pe3i L=3.5e-07 W=4.9e-06 AD=2.7195e-12 AS=2.7195e-12 PD=1.091e-05 PS=1.091e-05 $X=4595 $Y=186615 $dt=1
M26 18 EN VDD3I VDD3I pe3i L=3.5e-07 W=2.16e-06 AD=1.0368e-12 AS=1.0368e-12 PD=5.28e-06 PS=5.28e-06 $X=7005 $Y=254785 $dt=1
M27 22 14 VDDOI VDDOI pe3i L=3.5e-07 W=5e-06 AD=1.725e-12 AS=2.775e-12 PD=5.69e-06 PS=1.111e-05 $X=7245 $Y=186615 $dt=1
M28 VDDOI 14 22 VDDOI pe3i L=3.5e-07 W=5e-06 AD=1.725e-12 AS=1.725e-12 PD=5.69e-06 PS=5.69e-06 $X=8285 $Y=186615 $dt=1
M29 14 17 VDDOI VDDOI pe3i L=3.5e-07 W=2.6e-06 AD=7.02e-13 AS=1.248e-12 PD=3.14e-06 PS=6.16e-06 $X=8635 $Y=234395 $dt=1
M30 17 A VDD3I VDD3I pe3i L=3.5e-07 W=2.16e-06 AD=5.832e-13 AS=1.0368e-12 PD=2.7e-06 PS=5.28e-06 $X=8640 $Y=254785 $dt=1
M31 22 14 VDDOI VDDOI pe3i L=3.5e-07 W=5e-06 AD=1.725e-12 AS=1.725e-12 PD=5.69e-06 PS=5.69e-06 $X=9325 $Y=186615 $dt=1
M32 VDDOI 17 14 VDDOI pe3i L=3.5e-07 W=2.6e-06 AD=7.02e-13 AS=7.02e-13 PD=3.14e-06 PS=3.14e-06 $X=9525 $Y=234395 $dt=1
M33 VDD3I 18 17 VDD3I pe3i L=3.5e-07 W=2.16e-06 AD=1.0368e-12 AS=5.832e-13 PD=5.28e-06 PS=2.7e-06 $X=9530 $Y=254785 $dt=1
M34 VDDOI 14 22 VDDOI pe3i L=3.5e-07 W=5e-06 AD=2.775e-12 AS=1.725e-12 PD=1.111e-05 PS=5.69e-06 $X=10365 $Y=186615 $dt=1
M35 14 17 VDDOI VDDOI pe3i L=3.5e-07 W=2.6e-06 AD=7.02e-13 AS=7.02e-13 PD=3.14e-06 PS=3.14e-06 $X=10415 $Y=234395 $dt=1
M36 VDDOI 17 14 VDDOI pe3i L=3.5e-07 W=2.6e-06 AD=7.02e-13 AS=7.02e-13 PD=3.14e-06 PS=3.14e-06 $X=11305 $Y=234395 $dt=1
M37 16 20 VDDOI VDDOI pe3i L=3.5e-07 W=2.6e-06 AD=7.02e-13 AS=7.02e-13 PD=3.14e-06 PS=3.14e-06 $X=12195 $Y=234395 $dt=1
M38 VDDOI 20 16 VDDOI pe3i L=3.5e-07 W=2.6e-06 AD=7.02e-13 AS=7.02e-13 PD=3.14e-06 PS=3.14e-06 $X=13085 $Y=234395 $dt=1
M39 26 A VDD3I VDD3I pe3i L=3.5e-07 W=2.16e-06 AD=5.832e-13 AS=1.0368e-12 PD=2.7e-06 PS=5.28e-06 $X=13505 $Y=254785 $dt=1
M40 16 20 VDDOI VDDOI pe3i L=3.5e-07 W=2.6e-06 AD=7.02e-13 AS=7.02e-13 PD=3.14e-06 PS=3.14e-06 $X=13975 $Y=234395 $dt=1
M41 20 EN 26 VDD3I pe3i L=3.5e-07 W=2.16e-06 AD=1.0368e-12 AS=5.832e-13 PD=5.28e-06 PS=2.7e-06 $X=14395 $Y=254785 $dt=1
M42 VDDOI 20 16 VDDOI pe3i L=3.5e-07 W=2.6e-06 AD=1.248e-12 AS=7.02e-13 PD=6.16e-06 PS=3.14e-06 $X=14865 $Y=234395 $dt=1
M43 21 14 VDDOI VDDOI pe3i L=3.5e-07 W=5e-06 AD=1.725e-12 AS=2.775e-12 PD=5.69e-06 PS=1.111e-05 $X=59215 $Y=186615 $dt=1
M44 VDDOI 14 21 VDDOI pe3i L=3.5e-07 W=5e-06 AD=1.725e-12 AS=1.725e-12 PD=5.69e-06 PS=5.69e-06 $X=60255 $Y=186615 $dt=1
M45 21 14 VDDOI VDDOI pe3i L=3.5e-07 W=5e-06 AD=1.725e-12 AS=1.725e-12 PD=5.69e-06 PS=5.69e-06 $X=61295 $Y=186615 $dt=1
M46 VDDOI 14 21 VDDOI pe3i L=3.5e-07 W=5e-06 AD=2.775e-12 AS=1.725e-12 PD=1.111e-05 PS=5.69e-06 $X=62335 $Y=186615 $dt=1
M47 27 16 23 VDDOI pe3i L=4e-07 W=6.7e-06 AD=2.144e-12 AS=3.551e-12 PD=7.34e-06 PS=1.446e-05 $X=64050 $Y=186615 $dt=1
M48 VDDOI 16 27 VDDOI pe3i L=4e-07 W=6.7e-06 AD=3.551e-12 AS=2.144e-12 PD=1.446e-05 PS=7.34e-06 $X=65090 $Y=186615 $dt=1
R49 11 VDDOI L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=VDDOI $X=14380 $Y=198475 $dt=7
D50 11 VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=13360 $Y=198475 $dt=12
D51 VDDOI VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=17680 $Y=198475 $dt=12
.ends BT4PC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_pcutdio_pc                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_pcutdio_pc 1 2
** N=5 EP=2 FDC=2
D0 2 1 dp3 AREA=5.88986e-11 PJ=6.40282e-05 perimeter=6.40282e-05 $X=2765 $Y=76075 $dt=10
D1 1 2 dp3 AREA=5.88986e-11 PJ=6.40282e-05 perimeter=6.40282e-05 $X=37455 $Y=78455 $dt=10
.ends jio_pcutdio_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: PWRCUTDCPC                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt PWRCUTDCPC GNDOI1 PSUB GNDOI2 VDD3I1 VDDOI1 GNDI1 GNDI2 VDD3I2 VDDOI2 VDDRI1
+ GNDRI1 VDDRI2 GNDRI2
** N=20 EP=13 FDC=31
X80 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 0 0 0 $X=1370 $Y=75245
X81 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 4760 0 0 $X=1370 $Y=80005
X82 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 9520 0 0 $X=1370 $Y=84765
X83 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 14280 0 0 $X=1370 $Y=89525
X84 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 19040 0 0 $X=1370 $Y=94285
X85 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 23800 0 0 $X=1370 $Y=99045
X86 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 28560 0 0 $X=1370 $Y=103805
X87 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 33320 0 0 $X=1370 $Y=108565
X88 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 38080 0 0 $X=1370 $Y=113325
X89 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 42840 0 0 $X=1370 $Y=118085
X90 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 47600 0 0 $X=1370 $Y=122845
X91 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 52360 0 0 $X=1370 $Y=127605
X92 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 57120 0 0 $X=1370 $Y=132365
X93 GNDOI1 GNDOI2 jio_pcutdio_pc $T=0 61880 0 0 $X=1370 $Y=137125
D0 GNDOI2 GNDOI1 dp3 AREA=5.88986e-11 PJ=6.40282e-05 perimeter=6.40282e-05 $X=2765 $Y=142715 $dt=10
D1 PSUB GNDOI1 p_dnw3 AREA=2.32916e-09 PJ=0.00020788 perimeter=0.00020788 $X=1310 $Y=74975 $dt=13
D2 PSUB GNDOI2 p_dnw3 AREA=2.32916e-09 PJ=0.00020788 perimeter=0.00020788 $X=36000 $Y=74975 $dt=13
.ends PWRCUTDCPC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_ne3isbc_pc                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_ne3isbc_pc 2 3 5 6
*.DEVICECLIMB
** N=9 EP=4 FDC=3
R0 5 3 L=3.35e-06 W=3e-05 $[rdn3] $SUB=2 $X=955 $Y=1825 $dt=5
R1 3 6 L=3.35e-06 W=3e-05 $[rdn3] $SUB=2 $X=4960 $Y=1825 $dt=5
D2 2 3 dn3 AREA=1.98e-11 PJ=1.32e-06 perimeter=1.32e-06 $X=4300 $Y=1825 $dt=9
.ends jio_ne3isbc_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: jio_crnentr_pc                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt jio_crnentr_pc 1 2 3
** N=28 EP=3 FDC=66
X165 3 2 7 8 jio_ne3isbc_pc $T=207490 108730 0 180 $X=197170 $Y=74825
X166 3 2 5 6 jio_ne3isbc_pc $T=207490 142530 0 180 $X=197170 $Y=108625
X167 3 2 11 12 jio_ne3isbc_pc $T=216490 108730 0 180 $X=206170 $Y=74825
X168 3 2 9 10 jio_ne3isbc_pc $T=216490 142530 0 180 $X=206170 $Y=108625
X169 3 2 15 16 jio_ne3isbc_pc $T=225490 108730 0 180 $X=215170 $Y=74825
X170 3 2 13 14 jio_ne3isbc_pc $T=225490 142530 0 180 $X=215170 $Y=108625
X171 3 2 19 20 jio_ne3isbc_pc $T=226650 108730 1 0 $X=225590 $Y=74825
X172 3 2 17 18 jio_ne3isbc_pc $T=226650 142530 1 0 $X=225590 $Y=108625
X173 3 2 23 24 jio_ne3isbc_pc $T=235650 108730 1 0 $X=234590 $Y=74825
X174 3 2 21 22 jio_ne3isbc_pc $T=235650 142530 1 0 $X=234590 $Y=108625
X175 3 2 27 28 jio_ne3isbc_pc $T=244650 108730 1 0 $X=243590 $Y=74825
X176 3 2 25 26 jio_ne3isbc_pc $T=244650 142530 1 0 $X=243590 $Y=108625
M0 8 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.89e-11 PD=6.001e-05 PS=6.126e-05 $X=198780 $Y=76905 $dt=0
M1 6 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.89e-11 PD=6.001e-05 PS=6.126e-05 $X=198780 $Y=110705 $dt=0
M2 3 4 7 3 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=206540 $Y=76905 $dt=0
M3 3 4 5 3 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=206540 $Y=110705 $dt=0
M4 12 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=207780 $Y=76905 $dt=0
M5 10 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=207780 $Y=110705 $dt=0
M6 3 4 11 3 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=215540 $Y=76905 $dt=0
M7 3 4 9 3 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=215540 $Y=110705 $dt=0
M8 16 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=216780 $Y=76905 $dt=0
M9 14 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=216780 $Y=110705 $dt=0
M10 3 4 15 3 ne3i L=4e-07 W=3e-05 AD=3.39e-11 AS=1.5e-13 PD=3.226e-05 PS=6.001e-05 $X=224540 $Y=76905 $dt=0
M11 3 4 13 3 ne3i L=4e-07 W=3e-05 AD=3.39e-11 AS=1.5e-13 PD=3.226e-05 PS=6.001e-05 $X=224540 $Y=110705 $dt=0
M12 19 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=3.39e-11 PD=6.001e-05 PS=3.226e-05 $X=227200 $Y=76905 $dt=0
M13 17 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=3.39e-11 PD=6.001e-05 PS=3.226e-05 $X=227200 $Y=110705 $dt=0
M14 3 4 20 3 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=234960 $Y=76905 $dt=0
M15 3 4 18 3 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=234960 $Y=110705 $dt=0
M16 23 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=236200 $Y=76905 $dt=0
M17 21 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=236200 $Y=110705 $dt=0
M18 3 4 24 3 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=243960 $Y=76905 $dt=0
M19 3 4 22 3 ne3i L=4e-07 W=3e-05 AD=1.26e-11 AS=1.5e-13 PD=3.084e-05 PS=6.001e-05 $X=243960 $Y=110705 $dt=0
M20 27 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=245200 $Y=76905 $dt=0
M21 25 4 3 3 ne3i L=4e-07 W=3e-05 AD=1.5e-13 AS=1.26e-11 PD=6.001e-05 PS=3.084e-05 $X=245200 $Y=110705 $dt=0
M22 3 4 28 3 ne3i L=4e-07 W=3e-05 AD=1.89e-11 AS=1.5e-13 PD=6.126e-05 PS=6.001e-05 $X=252960 $Y=76905 $dt=0
M23 3 4 26 3 ne3i L=4e-07 W=3e-05 AD=1.89e-11 AS=1.5e-13 PD=6.126e-05 PS=6.001e-05 $X=252960 $Y=110705 $dt=0
D24 1 2 ddnwmv AREA=4.69976e-09 PJ=0.00027464 perimeter=0.00027464 $X=193640 $Y=72575 $dt=2
D25 3 2 dipdnwmv AREA=4.16648e-09 PJ=0.00025864 perimeter=0.00025864 $X=195640 $Y=74575 $dt=4
R26 4 3 L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=2 $X=256135 $Y=151635 $dt=6
D27 4 2 p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=256135 $Y=150615 $dt=11
D28 3 2 p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=256135 $Y=154935 $dt=11
D29 1 2 p_dnw3 AREA=1.44615e-11 PJ=1.709e-05 perimeter=1.709e-05 $X=255425 $Y=150175 $dt=13
.ends jio_crnentr_pc

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: CORNERESDPC                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt CORNERESDPC PSUB GNDOI VDDOI GNDI VDD3I GNDRI VDDRI
** N=9 EP=7 FDC=132
X432 PSUB VDDOI GNDOI jio_crnentr_pc $T=0 0 1 90 $X=72565 $Y=191090
X433 PSUB VDDOI GNDOI jio_crnentr_pc $T=0 0 0 0 $X=191090 $Y=72565
.ends CORNERESDPC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: APR00DPC                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt APR00DPC PSUB VDDOI PAD GNDOI VDD3I GNDI VDDRI GNDRI
** N=42 EP=8 FDC=149
X1073 VDDOI PAD 18 17 jio_pe3isb_pc $T=14365 150990 1 180 $X=6700 $Y=149060
X1074 VDDOI PAD 16 15 jio_pe3isb_pc $T=14365 184790 1 180 $X=6700 $Y=182860
X1075 VDDOI PAD 14 13 jio_pe3isb_pc $T=20965 150990 1 180 $X=13300 $Y=149060
X1076 VDDOI PAD 12 11 jio_pe3isb_pc $T=20965 184790 1 180 $X=13300 $Y=182860
X1077 VDDOI PAD 26 25 jio_pe3isb_pc $T=27565 150990 1 180 $X=19900 $Y=149060
X1078 VDDOI PAD 24 23 jio_pe3isb_pc $T=27565 184790 1 180 $X=19900 $Y=182860
X1079 VDDOI PAD 22 21 jio_pe3isb_pc $T=34165 150990 1 180 $X=26500 $Y=149060
X1080 VDDOI PAD 20 19 jio_pe3isb_pc $T=34165 184790 1 180 $X=26500 $Y=182860
X1081 VDDOI PAD 34 33 jio_pe3isb_pc $T=35835 150990 0 0 $X=35120 $Y=149060
X1082 VDDOI PAD 32 31 jio_pe3isb_pc $T=35835 184790 0 0 $X=35120 $Y=182860
X1083 VDDOI PAD 30 29 jio_pe3isb_pc $T=42435 150990 0 0 $X=41720 $Y=149060
X1084 VDDOI PAD 28 27 jio_pe3isb_pc $T=42435 184790 0 0 $X=41720 $Y=182860
X1085 VDDOI PAD 42 41 jio_pe3isb_pc $T=49035 150990 0 0 $X=48320 $Y=149060
X1086 VDDOI PAD 40 39 jio_pe3isb_pc $T=49035 184790 0 0 $X=48320 $Y=182860
X1087 VDDOI PAD 38 37 jio_pe3isb_pc $T=55635 150990 0 0 $X=54920 $Y=149060
X1088 VDDOI PAD 36 35 jio_pe3isb_pc $T=55635 184790 0 0 $X=54920 $Y=182860
X1277 VDDOI GNDOI 10 10 10 PAD PSUB jio_base_ntr_pc $T=0 0 0 0 $X=2560 $Y=72565
M0 18 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=8060 $Y=152815 $dt=1
M1 16 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=8060 $Y=186615 $dt=1
M2 VDDOI 9 17 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=13370 $Y=152815 $dt=1
M3 VDDOI 9 15 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=13370 $Y=186615 $dt=1
M4 14 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=14660 $Y=152815 $dt=1
M5 12 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=14660 $Y=186615 $dt=1
M6 VDDOI 9 13 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=19970 $Y=152815 $dt=1
M7 VDDOI 9 11 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=19970 $Y=186615 $dt=1
M8 26 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=21260 $Y=152815 $dt=1
M9 24 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=21260 $Y=186615 $dt=1
M10 VDDOI 9 25 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=26570 $Y=152815 $dt=1
M11 VDDOI 9 23 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=26570 $Y=186615 $dt=1
M12 22 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=27860 $Y=152815 $dt=1
M13 20 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=27860 $Y=186615 $dt=1
M14 VDDOI 9 21 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=33170 $Y=152815 $dt=1
M15 VDDOI 9 19 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=33170 $Y=186615 $dt=1
M16 33 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=36480 $Y=152815 $dt=1
M17 31 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=36480 $Y=186615 $dt=1
M18 VDDOI 9 34 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=41790 $Y=152815 $dt=1
M19 VDDOI 9 32 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=41790 $Y=186615 $dt=1
M20 29 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=43080 $Y=152815 $dt=1
M21 27 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=43080 $Y=186615 $dt=1
M22 VDDOI 9 30 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=48390 $Y=152815 $dt=1
M23 VDDOI 9 28 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=48390 $Y=186615 $dt=1
M24 41 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=49680 $Y=152815 $dt=1
M25 39 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=49680 $Y=186615 $dt=1
M26 VDDOI 9 42 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=54990 $Y=152815 $dt=1
M27 VDDOI 9 40 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=54990 $Y=186615 $dt=1
M28 37 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=56280 $Y=152815 $dt=1
M29 35 9 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=56280 $Y=186615 $dt=1
M30 VDDOI 9 38 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=61590 $Y=152815 $dt=1
M31 VDDOI 9 36 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=61590 $Y=186615 $dt=1
D32 PSUB VDDOI p_ddnwmv AREA=4.5084e-09 PJ=0.00026872 perimeter=0.00026872 $X=2500 $Y=150035 $dt=3
R33 9 VDDOI L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=VDDOI $X=4475 $Y=153720 $dt=7
R34 10 GNDOI L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=VDDOI $X=65085 $Y=153720 $dt=7
D35 9 VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=4475 $Y=152700 $dt=12
D36 VDDOI VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=4475 $Y=157020 $dt=12
D37 10 VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=65085 $Y=152700 $dt=12
D38 GNDOI VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=65085 $Y=157020 $dt=12
.ends APR00DPC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: APR04DPC                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt APR04DPC PSUB VDD3I VDDOI GNDOI GNDI PAD Y VDDRI GNDRI
** N=37 EP=9 FDC=139
X131 VDDOI PAD 17 16 jio_pe3isb_pc $T=14365 150990 1 180 $X=6700 $Y=149060
X132 VDDOI PAD 15 14 jio_pe3isb_pc $T=20965 150990 1 180 $X=13300 $Y=149060
X133 VDDOI PAD 25 24 jio_pe3isb_pc $T=27565 150990 1 180 $X=19900 $Y=149060
X134 VDDOI PAD 23 22 jio_pe3isb_pc $T=27565 184790 1 180 $X=19900 $Y=182860
X135 VDDOI PAD 21 20 jio_pe3isb_pc $T=34165 150990 1 180 $X=26500 $Y=149060
X136 VDDOI PAD 19 18 jio_pe3isb_pc $T=34165 184790 1 180 $X=26500 $Y=182860
X137 VDDOI PAD 33 32 jio_pe3isb_pc $T=35835 150990 0 0 $X=35120 $Y=149060
X138 VDDOI PAD 31 30 jio_pe3isb_pc $T=35835 184790 0 0 $X=35120 $Y=182860
X139 VDDOI PAD 29 28 jio_pe3isb_pc $T=42435 150990 0 0 $X=41720 $Y=149060
X140 VDDOI PAD 27 26 jio_pe3isb_pc $T=42435 184790 0 0 $X=41720 $Y=182860
X141 VDDOI PAD 37 36 jio_pe3isb_pc $T=49035 150990 0 0 $X=48320 $Y=149060
X142 VDDOI PAD 35 34 jio_pe3isb_pc $T=55635 150990 0 0 $X=54920 $Y=149060
X400 VDDOI GNDOI 11 11 11 PAD PSUB jio_base_ntr_pc $T=0 0 0 0 $X=2560 $Y=72565
M0 11 10 GNDOI GNDOI ne3i L=4e-07 W=1.2e-06 AD=6.36e-13 AS=6.36e-13 PD=3.46e-06 PS=3.46e-06 $X=10900 $Y=212165 $dt=0
M1 12 GNDOI GNDOI GNDOI ne3i L=4e-07 W=1.2e-05 AD=6e-14 AS=6.66e-12 PD=2.401e-05 PS=2.511e-05 $X=59470 $Y=203135 $dt=0
M2 GNDOI GNDOI 13 GNDOI ne3i L=4e-07 W=1.2e-05 AD=6.66e-12 AS=6e-14 PD=2.511e-05 PS=2.401e-05 $X=63170 $Y=203135 $dt=0
M3 17 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=8060 $Y=152815 $dt=1
M4 VDDOI 10 16 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=13370 $Y=152815 $dt=1
M5 15 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=14660 $Y=152815 $dt=1
M6 VDDOI 10 14 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=19970 $Y=152815 $dt=1
M7 25 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=21260 $Y=152815 $dt=1
M8 23 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=21260 $Y=186615 $dt=1
M9 VDDOI 10 24 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=26570 $Y=152815 $dt=1
M10 VDDOI 10 22 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=26570 $Y=186615 $dt=1
M11 21 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=27860 $Y=152815 $dt=1
M12 19 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=27860 $Y=186615 $dt=1
M13 VDDOI 10 20 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=33170 $Y=152815 $dt=1
M14 VDDOI 10 18 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=33170 $Y=186615 $dt=1
M15 32 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=36480 $Y=152815 $dt=1
M16 30 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=2.04e-11 PD=6.001e-05 PS=6.136e-05 $X=36480 $Y=186615 $dt=1
M17 VDDOI 10 33 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=41790 $Y=152815 $dt=1
M18 VDDOI 10 31 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=41790 $Y=186615 $dt=1
M19 28 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=43080 $Y=152815 $dt=1
M20 26 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=43080 $Y=186615 $dt=1
M21 VDDOI 10 29 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=48390 $Y=152815 $dt=1
M22 VDDOI 10 27 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=48390 $Y=186615 $dt=1
M23 36 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=49680 $Y=152815 $dt=1
M24 Y VDDOI VDDOI VDDOI pe3i L=3.5e-07 W=1.2e-05 AD=6.78e-12 AS=6.24e-12 PD=1.313e-05 PS=2.504e-05 $X=51820 $Y=202785 $dt=1
M25 VDDOI VDDOI Y VDDOI pe3i L=3.5e-07 W=1.2e-05 AD=6.24e-12 AS=6.78e-12 PD=2.504e-05 PS=1.313e-05 $X=53300 $Y=202785 $dt=1
M26 VDDOI 10 37 VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.41e-11 AS=1.5e-13 PD=3.094e-05 PS=6.001e-05 $X=54990 $Y=152815 $dt=1
M27 34 10 VDDOI VDDOI pe3i L=3.5e-07 W=3e-05 AD=1.5e-13 AS=1.41e-11 PD=6.001e-05 PS=3.094e-05 $X=56280 $Y=152815 $dt=1
M28 VDDOI 10 35 VDDOI pe3i L=3.5e-07 W=3e-05 AD=2.04e-11 AS=1.5e-13 PD=6.136e-05 PS=6.001e-05 $X=61590 $Y=152815 $dt=1
D29 PSUB VDDOI ddnwmv AREA=9.8345e-10 PJ=0.00016026 perimeter=0.00016026 $X=2500 $Y=224395 $dt=2
D30 PSUB VDD3I ddnwmv AREA=9.789e-10 PJ=0.00016012 perimeter=0.00016012 $X=2500 $Y=244525 $dt=2
D31 PSUB VDDOI p_ddnwmv AREA=4.5084e-09 PJ=0.00026872 perimeter=0.00026872 $X=2500 $Y=150035 $dt=3
D32 GNDOI VDDOI dipdnwmv AREA=2.1664e-10 PJ=5.908e-05 perimeter=5.908e-05 $X=4500 $Y=201395 $dt=4
D33 GNDOI VDDOI dipdnwmv AREA=1.2696e-10 PJ=4.787e-05 perimeter=4.787e-05 $X=57565 $Y=201395 $dt=4
R34 12 Y L=1.32e-06 W=1.2e-05 $[rdn3] $SUB=GNDOI $X=59875 $Y=203135 $dt=5
R35 Y 13 L=1.32e-06 W=1.2e-05 $[rdn3] $SUB=GNDOI $X=61850 $Y=203135 $dt=5
R36 10 VDDOI L=3.3e-06 W=4.4e-07 $[rdp3] $SUB=VDDOI $X=14380 $Y=198475 $dt=7
D37 GNDOI Y dn3 AREA=7.92e-12 PJ=1.32e-06 perimeter=1.32e-06 $X=61190 $Y=203135 $dt=9
D38 10 VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=13360 $Y=198475 $dt=12
D39 VDDOI VDDOI p_dp3 AREA=4.488e-13 PJ=2.48e-06 perimeter=2.48e-06 $X=17680 $Y=198475 $dt=12
R40 PAD Y L=2.2e-06 W=2e-06 $[rpp1] $X=60020 $Y=189980 $dt=14
.ends APR04DPC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ioring3                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ioring3 CLK ENABLE GNDA GNDD GNDOR GNDORA INL OUT0 OUT1 OUT2
+ OUTL PSUB RESET VDDA VDDD VDDOR VDDORA clk_core enable_core inl_core
+ out0_core out1_core out2_core reset_core
** N=38 EP=24 FDC=2805
X8 PSUB GNDOR VDDOR VDDD GNDD VDDOR GNDOR PSUBPADPC $T=352460 40295 0 0 $X=352140 $Y=40295
X9 VDDD GNDD VDDOR VDDOR GNDOR GNDOR PSUB VDDPADPC $T=282460 40295 0 0 $X=282140 $Y=40295
X10 VDDA GNDA VDDORA VDDORA GNDORA GNDORA PSUB VDDPADPC $T=1122460 40295 0 0 $X=1122140 $Y=40295
X11 PSUB VDDOR GNDOR VDDD GNDD GNDOR VDDORPADPC $T=212460 40295 0 0 $X=212140 $Y=40295
X12 PSUB VDDORA GNDORA VDDA GNDA GNDORA VDDORPADPC $T=1052460 40295 0 0 $X=1052140 $Y=40295
X13 GNDD VDDD VDDOR VDDOR GNDOR GNDOR PSUB GNDPADPC $T=72460 40295 0 0 $X=72140 $Y=40295
X14 GNDA VDDA VDDORA VDDORA GNDORA GNDORA PSUB GNDPADPC $T=982460 40295 0 0 $X=982140 $Y=40295
X15 PSUB VDDOR GNDOR VDDD GNDD VDDOR GNDORPADPC $T=142460 40295 0 0 $X=142140 $Y=40295
X16 PSUB VDDORA GNDORA VDDA GNDA VDDORA GNDORPADPC $T=912460 40295 0 0 $X=912140 $Y=40295
X17 VDDOR VDDD PSUB GNDD GNDOR VDDOR GNDOR enable_core ENABLE 13
+ GNDD ICPC $T=422460 40295 0 0 $X=422140 $Y=40295
X18 VDDOR VDDD PSUB GNDD GNDOR VDDOR GNDOR clk_core CLK 16
+ GNDD ICPC $T=492460 40295 0 0 $X=492140 $Y=40295
X19 VDDOR VDDD PSUB GNDD GNDOR VDDOR GNDOR reset_core RESET 19
+ GNDD ICPC $T=562460 40295 0 0 $X=562140 $Y=40295
X20 VDDD VDDOR GNDOR out0_core PSUB GNDD GNDD VDDOR GNDOR OUT0 BT4PC $T=632460 40295 0 0 $X=632140 $Y=40295
X21 VDDD VDDOR GNDOR out1_core PSUB GNDD GNDD VDDOR GNDOR OUT1 BT4PC $T=702460 40295 0 0 $X=702140 $Y=40295
X22 VDDD VDDOR GNDOR out2_core PSUB GNDD GNDD VDDOR GNDOR OUT2 BT4PC $T=772460 40295 0 0 $X=772140 $Y=40295
X23 2 PSUB GNDOR 26 27 28 GNDD VDDD VDDOR 29
+ 30 VDDOR GNDOR PWRCUTDCPC $T=-258540 371295 0 270 $X=-187155 $Y=300975
X24 GNDOR PSUB GNDORA VDDD VDDOR GNDD GNDA VDDA VDDORA VDDOR
+ GNDOR VDDORA GNDORA PWRCUTDCPC $T=842460 40295 0 0 $X=842140 $Y=111680
X25 GNDORA PSUB 2 VDDA VDDORA GNDA 31 32 33 VDDORA
+ GNDORA 34 35 PWRCUTDCPC $T=1663460 301295 0 90 $X=1402140 $Y=300975
X28 PSUB GNDOR VDDOR GNDD VDDD GNDOR VDDOR CORNERESDPC $T=-258540 40295 0 0 $X=-187155 $Y=111680
X29 PSUB GNDORA VDDORA GNDA VDDA GNDORA VDDORA CORNERESDPC $T=1663460 40295 0 90 $X=1402140 $Y=111680
X30 PSUB VDDORA OUTL GNDORA VDDA GNDA VDDORA GNDORA APR00DPC $T=1262460 40295 0 0 $X=1262140 $Y=40295
X31 PSUB VDDA VDDORA GNDORA GNDA INL inl_core VDDORA GNDORA APR04DPC $T=1192460 40295 0 0 $X=1192140 $Y=40295
.ends ioring3
